* NGSPICE file created from divider.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt divider A[0] A[10] A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19] A[1]
+ A[20] A[21] A[22] A[23] A[24] A[25] A[26] A[27] A[28] A[29] A[2] A[30] A[31] A[3]
+ A[4] A[5] A[6] A[7] A[8] A[9] B[0] B[10] B[11] B[12] B[13] B[14] B[15] B[16] B[17]
+ B[18] B[19] B[1] B[20] B[21] B[22] B[23] B[24] B[25] B[26] B[27] B[28] B[29] B[2]
+ B[30] B[31] B[3] B[4] B[5] B[6] B[7] B[8] B[9] D[0] D[10] D[11] D[12] D[13] D[14]
+ D[15] D[16] D[17] D[18] D[19] D[1] D[20] D[21] D[22] D[23] D[24] D[25] D[26] D[27]
+ D[28] D[29] D[2] D[30] D[31] D[3] D[4] D[5] D[6] D[7] D[8] D[9] R[0] R[10] R[11]
+ R[12] R[13] R[14] R[15] R[16] R[17] R[18] R[19] R[1] R[20] R[21] R[22] R[23] R[24]
+ R[25] R[26] R[27] R[28] R[29] R[2] R[30] R[31] R[3] R[4] R[5] R[6] R[7] R[8] R[9]
+ VGND VPWR clk err ok reset start
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1270_ clknet_3_5__leaf_clk _0108_ _0012_ VGND VGND VPWR VPWR reg32_denom.bit6.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0985_ _0461_ VGND VGND VPWR VPWR reg32_result.bit14.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0770_ _0205_ _0203_ _0292_ _0202_ _0212_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1322_ clknet_3_2__leaf_clk reg32_work.bit27.BitData _0064_ VGND VGND VPWR VPWR net118
+ sky130_fd_sc_hd__dfrtp_4
X_1253_ _0151_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_1184_ _0563_ _0564_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and2b_1
X_0968_ _0452_ VGND VGND VPWR VPWR reg32_result.bit6.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ _0216_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ reg32_denom.bit3.BitOut net121 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__and2b_1
X_0753_ _0268_ _0271_ _0272_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o21ai_1
X_0684_ _0205_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ clknet_3_5__leaf_clk reg32_work.bit10.BitData _0047_ VGND VGND VPWR VPWR net100
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1236_ _0140_ _0141_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1098_ _0515_ _0516_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__and2b_1
X_1167_ _0491_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ net39 net38 net37 net36 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or4_1
X_0805_ reg32_denom.bit31.BitOut _0324_ _0323_ _0326_ _0327_ VGND VGND VPWR VPWR _0328_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0667_ net136 net137 _0193_ VGND VGND VPWR VPWR cycle_reg.bit1.BitData sky130_fd_sc_hd__a21o_1
X_0598_ net58 reg32_denom.bit3.BitOut _0154_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
X_0736_ reg32_denom.bit12.BitOut net101 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nor2b_1
X_1219_ _0592_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 reg32_denom.bit5.BitOut VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ net17 net82 _0191_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0719_ net126 reg32_denom.bit6.BitOut VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput75 net75 VGND VGND VPWR VPWR D[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput97 net97 VGND VGND VPWR VPWR D[8] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR D[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0984_ net6 net149 _0459_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1321_ clknet_3_2__leaf_clk reg32_work.bit26.BitData _0063_ VGND VGND VPWR VPWR net117
+ sky130_fd_sc_hd__dfrtp_2
X_1252_ _0140_ _0141_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__and2b_1
X_1183_ _0572_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0967_ net29 net94 _0448_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux2_1
X_0898_ reg32_denom.bit18.BitOut _0289_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o21ba_1
X_0752_ net100 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__inv_2
X_0821_ _0229_ _0233_ _0227_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o21ai_1
X_0683_ net109 reg32_denom.bit20.BitOut VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2b_1
X_1304_ clknet_3_7__leaf_clk reg32_work.bit9.BitData _0046_ VGND VGND VPWR VPWR net130
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1235_ _0142_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_1166_ _0489_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__buf_2
X_1097_ _0525_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ net35 net34 net44 net63 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or4_1
X_0735_ _0256_ _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__nand2_1
X_0804_ reg32_denom.bit31.BitOut _0324_ _0319_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21bo_1
X_0597_ _0156_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
X_0666_ cycle_reg.bit0.BitOut cycle_reg.bit1.BitOut _0192_ VGND VGND VPWR VPWR _0193_
+ sky130_fd_sc_hd__o21ai_1
X_1218_ _0587_ _0588_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2b_1
X_1149_ _0554_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold31 reg32_denom.bit26.BitOut VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net105 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1003_ _0470_ VGND VGND VPWR VPWR reg32_result.bit23.BitData sky130_fd_sc_hd__clkbuf_1
X_0718_ reg32_denom.bit6.BitOut net126 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0649_ net60 net163 _0182_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
Xoutput76 net76 VGND VGND VPWR VPWR D[18] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR D[28] sky130_fd_sc_hd__buf_2
Xoutput98 net98 VGND VGND VPWR VPWR D[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0983_ _0460_ VGND VGND VPWR VPWR reg32_result.bit13.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ clknet_3_2__leaf_clk reg32_work.bit25.BitData _0062_ VGND VGND VPWR VPWR net116
+ sky130_fd_sc_hd__dfrtp_2
X_1182_ _0563_ _0564_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and2b_1
X_1251_ _0150_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0966_ _0451_ VGND VGND VPWR VPWR reg32_result.bit5.BitData sky130_fd_sc_hd__clkbuf_1
X_0897_ _0398_ _0217_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0751_ _0267_ _0270_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0820_ net148 _0337_ _0340_ _0190_ VGND VGND VPWR VPWR reg32_work.bit2.BitData sky130_fd_sc_hd__o211a_1
X_1303_ clknet_3_7__leaf_clk reg32_work.bit8.BitData _0045_ VGND VGND VPWR VPWR net129
+ sky130_fd_sc_hd__dfrtp_1
X_0682_ reg32_denom.bit20.BitOut net109 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2b_2
X_1096_ _0515_ _0516_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__and2b_1
X_1165_ _0562_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_1234_ _0140_ _0141_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__and2b_1
X_0949_ _0440_ _0441_ _0347_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0803_ _0315_ _0325_ _0314_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a21o_1
X_0665_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0734_ reg32_denom.bit13.BitOut net102 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or2b_1
X_0596_ net56 reg32_denom.bit30.BitOut _0154_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
X_1217_ _0591_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_1148_ _0551_ _0552_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2b_1
X_1079_ _0491_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__buf_2
Xhold32 net78 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net106 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 reg32_denom.bit1.BitOut VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1002_ net16 net81 _0191_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0648_ _0183_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
X_0717_ _0236_ _0239_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR D[19] sky130_fd_sc_hd__clkbuf_4
Xoutput88 net88 VGND VGND VPWR VPWR D[29] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 VGND VGND VPWR VPWR R[0] sky130_fd_sc_hd__clkbuf_4
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0982_ net5 net70 _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1250_ _0140_ _0141_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__and2b_1
X_1181_ _0571_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0896_ net132 _0400_ VGND VGND VPWR VPWR reg32_work.bit18.BitData sky130_fd_sc_hd__nor2_1
X_0965_ net28 net93 _0448_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0750_ _0271_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0681_ _0202_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2b_1
X_1302_ clknet_3_5__leaf_clk reg32_work.bit7.BitData _0044_ VGND VGND VPWR VPWR net128
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1233_ net66 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1095_ _0524_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_1164_ _0551_ _0552_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and2b_1
X_0948_ _0318_ _0326_ _0321_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a21oi_2
X_0879_ reg32_denom.bit14.BitOut net103 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0802_ reg32_denom.bit28.BitOut net118 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or2b_1
X_0733_ net102 reg32_denom.bit13.BitOut VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0664_ u1.q VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_4
X_1216_ _0587_ _0588_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0595_ _0155_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
X_1147_ _0553_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
X_1078_ _0489_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 net129 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 reg32_denom.bit27.BitOut VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 reg32_denom.bit20.BitOut VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
X_1001_ _0469_ VGND VGND VPWR VPWR reg32_result.bit22.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0647_ net61 net160 _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
X_0716_ _0237_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput67 net67 VGND VGND VPWR VPWR D[0] sky130_fd_sc_hd__clkbuf_4
Xoutput78 net78 VGND VGND VPWR VPWR D[1] sky130_fd_sc_hd__buf_2
Xoutput89 net89 VGND VGND VPWR VPWR D[2] sky130_fd_sc_hd__clkbuf_4
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0981_ u1.q VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1180_ _0563_ _0564_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0964_ _0450_ VGND VGND VPWR VPWR reg32_result.bit4.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0895_ _0289_ _0399_ _0329_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0680_ reg32_denom.bit21.BitOut net111 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__or2b_1
X_1301_ clknet_3_5__leaf_clk reg32_work.bit6.BitData _0043_ VGND VGND VPWR VPWR net127
+ sky130_fd_sc_hd__dfrtp_4
X_1232_ net65 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1094_ _0515_ _0516_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__and2b_1
X_1163_ _0561_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0947_ _0318_ _0321_ _0326_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0878_ _0386_ VGND VGND VPWR VPWR reg32_work.bit14.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0801_ net122 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__inv_2
X_0594_ net64 reg32_denom.bit9.BitOut _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
X_0663_ u1.q VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__inv_2
X_0732_ reg32_denom.bit15.BitOut net104 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__xor2_2
X_1215_ _0590_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_1146_ _0551_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__and2b_1
X_1077_ _0514_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 net120 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 reg32_denom.bit0.BitOut VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
X_1000_ net15 net80 _0459_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
X_0715_ net124 reg32_denom.bit4.BitOut VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__and2b_1
X_0646_ u1.q VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__buf_4
X_1129_ _0543_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput68 net68 VGND VGND VPWR VPWR D[10] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR D[20] sky130_fd_sc_hd__buf_2
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0629_ _0173_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0980_ _0458_ VGND VGND VPWR VPWR reg32_result.bit12.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0894_ _0217_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__xor2_1
X_0963_ net27 net92 _0448_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _0139_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_1300_ clknet_3_5__leaf_clk reg32_work.bit5.BitData _0042_ VGND VGND VPWR VPWR net126
+ sky130_fd_sc_hd__dfrtp_2
X_1162_ _0551_ _0552_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__and2b_1
X_1093_ _0523_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
X_0946_ net119 _0338_ _0437_ _0439_ _0192_ VGND VGND VPWR VPWR reg32_work.bit29.BitData
+ sky130_fd_sc_hd__o221a_1
X_0877_ _0192_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0800_ _0321_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0731_ reg32_denom.bit14.BitOut net103 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__xor2_2
X_0593_ u1.q VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_4
X_0662_ _0190_ net136 VGND VGND VPWR VPWR cycle_reg.bit0.BitData sky130_fd_sc_hd__nand2_1
X_1214_ _0587_ _0588_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__and2b_1
X_1145_ _0491_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__buf_2
X_1076_ _0503_ _0504_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__and2b_1
X_0929_ net115 _0394_ _0426_ _0391_ VGND VGND VPWR VPWR reg32_work.bit25.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 net114 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0331_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0714_ reg32_denom.bit4.BitOut net124 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__and2b_1
X_0645_ _0181_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_1128_ _0539_ _0540_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2b_1
X_1059_ _0505_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput69 net69 VGND VGND VPWR VPWR D[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0628_ net39 reg32_denom.bit15.BitOut _0171_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0962_ _0449_ VGND VGND VPWR VPWR reg32_result.bit3.BitData sky130_fd_sc_hd__clkbuf_1
X_0893_ _0221_ _0224_ _0286_ _0288_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _0587_ _0588_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__and2b_1
X_1092_ _0515_ _0516_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and2b_1
X_1161_ _0560_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0945_ _0347_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nand2_1
X_0876_ net103 _0384_ net133 VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1359_ clknet_3_3__leaf_clk reg32_result.bit31.BitData _0101_ VGND VGND VPWR VPWR
+ net91 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0730_ _0240_ _0248_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a21oi_2
X_0661_ _0154_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_4
X_1213_ _0589_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
X_1144_ _0489_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__buf_2
X_1075_ _0513_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
X_0859_ _0266_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__inv_2
X_0928_ _0347_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nand2_1
Xhold14 net72 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 reg32_work.bit0.BitData VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0644_ net62 reg32_denom.bit7.BitOut _0171_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
X_0713_ _0226_ _0229_ _0233_ _0234_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o311ai_2
X_1127_ _0542_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
X_1058_ _0503_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0627_ _0172_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0961_ net26 net152 _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0892_ net143 _0394_ _0397_ _0391_ VGND VGND VPWR VPWR reg32_work.bit17.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1160_ _0551_ _0552_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and2b_1
X_1091_ _0522_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_0944_ _0325_ _0434_ _0316_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21o_1
X_0875_ _0254_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__xor2_1
X_1358_ clknet_3_3__leaf_clk reg32_result.bit30.BitData _0100_ VGND VGND VPWR VPWR
+ net90 sky130_fd_sc_hd__dfrtp_1
X_1289_ clknet_3_0__leaf_clk _0127_ _0031_ VGND VGND VPWR VPWR reg32_denom.bit25.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_0660_ _0189_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_1212_ _0587_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__and2b_1
X_1143_ _0550_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
X_1074_ _0503_ _0504_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0927_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0858_ _0370_ VGND VGND VPWR VPWR reg32_work.bit10.BitData sky130_fd_sc_hd__clkbuf_1
X_0789_ _0297_ _0299_ _0303_ _0311_ _0296_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a221o_1
Xhold26 reg32_denom.bit24.BitOut VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net110 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0712_ reg32_denom.bit3.BitOut net121 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or2b_1
X_0643_ _0180_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
X_1126_ _0539_ _0540_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__and2b_1
X_1057_ _0491_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0626_ net40 reg32_denom.bit16.BitOut _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
X_1109_ _0532_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0609_ net49 net159 _0160_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0960_ u1.q VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0891_ _0347_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nand2_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _0515_ _0516_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0943_ _0316_ _0325_ _0434_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0874_ _0281_ _0259_ _0378_ _0256_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1288_ clknet_3_0__leaf_clk _0126_ _0030_ VGND VGND VPWR VPWR reg32_denom.bit24.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1357_ clknet_3_3__leaf_clk reg32_result.bit29.BitData _0099_ VGND VGND VPWR VPWR
+ net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1211_ net66 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__buf_2
X_1142_ _0539_ _0540_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and2b_1
X_1073_ _0512_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0857_ _0192_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__and2_1
X_0926_ _0304_ _0420_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold16 net71 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 reg32_denom.bit6.BitOut VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _0304_ _0310_ _0308_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0711_ reg32_denom.bit2.BitOut _0226_ net110 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0642_ net63 reg32_denom.bit8.BitOut _0171_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
X_1125_ _0541_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_1056_ _0489_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0909_ _0347_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0625_ u1.q VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1108_ _0527_ _0528_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2b_1
X_1039_ _0494_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0608_ _0162_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0890_ _0224_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ net138 _0394_ _0436_ _0391_ VGND VGND VPWR VPWR reg32_work.bit28.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_27_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0873_ _0338_ _0380_ _0381_ _0382_ VGND VGND VPWR VPWR reg32_work.bit13.BitData sky130_fd_sc_hd__a31oi_1
X_1287_ clknet_3_0__leaf_clk _0125_ _0029_ VGND VGND VPWR VPWR reg32_denom.bit23.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1356_ clknet_3_2__leaf_clk reg32_result.bit28.BitData _0098_ VGND VGND VPWR VPWR
+ net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1210_ net65 VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__clkbuf_2
X_1141_ _0549_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_1072_ _0503_ _0504_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0856_ net130 _0368_ net133 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
X_0787_ reg32_denom.bit25.BitOut net115 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__and2b_1
X_0925_ _0307_ _0308_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__nand2_1
Xhold28 net69 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 net121 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ clknet_3_7__leaf_clk reg32_result.bit11.BitData _0081_ VGND VGND VPWR VPWR
+ net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0710_ _0230_ _0231_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a21oi_2
X_0641_ _0179_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and2b_1
X_1055_ _0502_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0839_ _0192_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__and2_1
X_0908_ _0204_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0624_ _0170_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1107_ _0531_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1038_ _0490_ _0492_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0607_ net50 reg32_denom.bit25.BitOut _0160_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0941_ _0434_ _0435_ _0330_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0872_ net102 _0330_ _0192_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21ai_1
X_1355_ clknet_3_3__leaf_clk reg32_result.bit27.BitData _0097_ VGND VGND VPWR VPWR
+ net86 sky130_fd_sc_hd__dfrtp_2
X_1286_ clknet_3_0__leaf_clk _0124_ _0028_ VGND VGND VPWR VPWR reg32_denom.bit22.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ _0539_ _0540_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__and2b_1
X_1071_ _0511_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
X_0924_ net146 _0394_ _0422_ _0391_ VGND VGND VPWR VPWR reg32_work.bit24.BitData sky130_fd_sc_hd__o211a_1
X_0855_ _0266_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__xnor2_1
X_0786_ _0303_ _0306_ _0307_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1338_ clknet_3_7__leaf_clk reg32_result.bit10.BitData _0080_ VGND VGND VPWR VPWR
+ net68 sky130_fd_sc_hd__dfrtp_1
Xhold29 net108 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 net84 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ clknet_3_5__leaf_clk _0107_ _0011_ VGND VGND VPWR VPWR reg32_denom.bit5.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0640_ net44 net154 _0171_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
X_1123_ _0491_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__clkbuf_2
X_1054_ _0490_ _0492_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0907_ _0205_ _0406_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nand2_1
X_0838_ net126 _0354_ net133 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
X_0769_ _0291_ _0207_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0623_ net41 reg32_denom.bit17.BitOut _0160_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
X_1106_ _0527_ _0528_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1037_ _0493_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0606_ _0161_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0313_ _0317_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ _0258_ _0259_ _0378_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__or3_1
X_1285_ clknet_3_0__leaf_clk _0123_ _0027_ VGND VGND VPWR VPWR reg32_denom.bit21.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1354_ clknet_3_6__leaf_clk reg32_result.bit26.BitData _0096_ VGND VGND VPWR VPWR
+ net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ _0503_ _0504_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__and2b_1
X_0854_ _0268_ _0271_ _0360_ _0272_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o31a_1
X_0923_ _0420_ _0421_ _0347_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o21ai_1
X_0785_ net115 reg32_denom.bit25.BitOut VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1268_ clknet_3_4__leaf_clk _0106_ _0010_ VGND VGND VPWR VPWR reg32_denom.bit4.BitOut
+ sky130_fd_sc_hd__dfrtp_1
Xhold19 net89 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ clknet_3_3__leaf_clk reg32_result.bit9.BitData _0079_ VGND VGND VPWR VPWR
+ net98 sky130_fd_sc_hd__dfrtp_1
X_1199_ _0581_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1122_ _0489_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__clkbuf_2
X_1053_ _0501_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0837_ _0243_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0906_ net109 _0394_ _0408_ _0391_ VGND VGND VPWR VPWR reg32_work.bit20.BitData sky130_fd_sc_hd__o211a_1
X_0768_ reg32_denom.bit19.BitOut _0287_ _0288_ _0218_ _0290_ VGND VGND VPWR VPWR _0291_
+ sky130_fd_sc_hd__o221a_1
X_0699_ net106 reg32_denom.bit17.BitOut VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0622_ _0169_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
X_1105_ _0530_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_1036_ _0490_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0605_ net51 net164 _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
X_1019_ _0478_ VGND VGND VPWR VPWR reg32_result.bit31.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0870_ _0259_ _0378_ _0258_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__o21ai_1
X_1284_ clknet_3_0__leaf_clk _0122_ _0026_ VGND VGND VPWR VPWR reg32_denom.bit20.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1353_ clknet_3_6__leaf_clk reg32_result.bit25.BitData _0095_ VGND VGND VPWR VPWR
+ net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _0468_ VGND VGND VPWR VPWR reg32_result.bit21.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0853_ net144 _0337_ _0366_ _0190_ VGND VGND VPWR VPWR reg32_work.bit9.BitData sky130_fd_sc_hd__o211a_1
X_0922_ _0295_ _0306_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0784_ reg32_denom.bit25.BitOut net115 VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or2b_1
Xinput1 A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_1198_ _0575_ _0576_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__and2b_1
X_1336_ clknet_3_3__leaf_clk reg32_result.bit8.BitData _0078_ VGND VGND VPWR VPWR
+ net97 sky130_fd_sc_hd__dfrtp_1
X_1267_ clknet_3_1__leaf_clk _0105_ _0009_ VGND VGND VPWR VPWR reg32_denom.bit31.BitOut
+ sky130_fd_sc_hd__dfrtp_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1121_ _0538_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_1052_ _0490_ _0492_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0836_ _0237_ _0240_ _0246_ _0245_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ _0406_ _0407_ _0330_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0767_ reg32_denom.bit19.BitOut _0287_ _0289_ reg32_denom.bit18.BitOut VGND VGND
+ VPWR VPWR _0290_ sky130_fd_sc_hd__a211o_1
X_0698_ _0219_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ clknet_3_2__leaf_clk reg32_work.bit24.BitData _0061_ VGND VGND VPWR VPWR net115
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0621_ net42 reg32_denom.bit18.BitOut _0160_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1104_ _0527_ _0528_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1035_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0819_ _0338_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nand2_1
X_0604_ u1.q VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__buf_4
X_1018_ net25 net90 _0191_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1283_ clknet_3_1__leaf_clk _0121_ _0025_ VGND VGND VPWR VPWR reg32_denom.bit2.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1352_ clknet_3_6__leaf_clk reg32_result.bit24.BitData _0094_ VGND VGND VPWR VPWR
+ net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0998_ net14 net79 _0459_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0921_ _0295_ _0306_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and2_1
X_0852_ _0338_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nand2_1
X_0783_ _0304_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1335_ clknet_3_3__leaf_clk reg32_result.bit7.BitData _0077_ VGND VGND VPWR VPWR
+ net96 sky130_fd_sc_hd__dfrtp_2
Xinput2 A[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1197_ _0580_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_1266_ clknet_3_4__leaf_clk _0104_ _0008_ VGND VGND VPWR VPWR reg32_denom.bit29.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1051_ _0500_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
X_1120_ _0527_ _0528_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0904_ _0291_ _0207_ _0405_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0835_ net125 _0337_ _0352_ _0190_ VGND VGND VPWR VPWR reg32_work.bit5.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0766_ net107 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__inv_2
X_0697_ net105 reg32_denom.bit16.BitOut VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1318_ clknet_3_0__leaf_clk reg32_work.bit23.BitData _0060_ VGND VGND VPWR VPWR net114
+ sky130_fd_sc_hd__dfrtp_1
X_1249_ _0149_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0620_ _0168_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_1034_ net66 VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__buf_2
X_1103_ _0529_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput60 B[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlymetal6s2s_1
X_0749_ net129 reg32_denom.bit9.BitOut VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0818_ _0229_ _0233_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0603_ _0159_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1017_ _0477_ VGND VGND VPWR VPWR reg32_result.bit30.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1351_ clknet_3_3__leaf_clk reg32_result.bit23.BitData _0093_ VGND VGND VPWR VPWR
+ net82 sky130_fd_sc_hd__dfrtp_2
X_1282_ clknet_3_1__leaf_clk _0120_ _0024_ VGND VGND VPWR VPWR reg32_denom.bit18.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0997_ _0467_ VGND VGND VPWR VPWR reg32_result.bit20.BitData sky130_fd_sc_hd__clkbuf_1
X_0920_ net113 _0394_ _0417_ _0419_ _0192_ VGND VGND VPWR VPWR reg32_work.bit23.BitData
+ sky130_fd_sc_hd__o221a_1
X_0851_ _0273_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__xnor2_1
X_0782_ net114 reg32_denom.bit24.BitOut VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1334_ clknet_3_2__leaf_clk reg32_result.bit6.BitData _0076_ VGND VGND VPWR VPWR
+ net95 sky130_fd_sc_hd__dfrtp_1
X_1265_ clknet_3_1__leaf_clk _0103_ _0007_ VGND VGND VPWR VPWR reg32_denom.bit19.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1196_ _0575_ _0576_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__and2b_1
Xinput3 A[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1050_ _0490_ _0492_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0834_ _0338_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nand2_1
X_0903_ _0291_ _0405_ _0207_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0765_ _0223_ _0219_ _0222_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21bo_1
X_0696_ reg32_denom.bit16.BitOut net105 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__or2b_1
X_1317_ clknet_3_1__leaf_clk reg32_work.bit22.BitData _0059_ VGND VGND VPWR VPWR net113
+ sky130_fd_sc_hd__dfrtp_2
X_1248_ _0140_ _0141_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__and2b_1
X_1179_ _0570_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ _0527_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1033_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__buf_2
Xinput50 B[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 B[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XFILLER_0_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0817_ _0330_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_4
X_0748_ reg32_denom.bit9.BitOut net129 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__and2b_1
X_0679_ net111 reg32_denom.bit21.BitOut VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0602_ net52 net155 _0154_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1016_ net24 net88 _0191_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1281_ clknet_3_1__leaf_clk _0119_ _0023_ VGND VGND VPWR VPWR reg32_denom.bit17.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1350_ clknet_3_3__leaf_clk reg32_result.bit22.BitData _0092_ VGND VGND VPWR VPWR
+ net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ net13 net77 _0459_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0850_ _0268_ _0360_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__nor2_1
X_0781_ reg32_denom.bit24.BitOut net114 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 A[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_1333_ clknet_3_2__leaf_clk reg32_result.bit5.BitData _0075_ VGND VGND VPWR VPWR
+ net94 sky130_fd_sc_hd__dfrtp_1
X_1264_ clknet_3_4__leaf_clk _0102_ _0006_ VGND VGND VPWR VPWR reg32_denom.bit0.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1195_ _0579_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0979_ net4 net161 _0448_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0833_ _0349_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__xnor2_1
X_0902_ _0225_ _0286_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or2_1
X_0764_ net108 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__inv_2
X_0695_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1316_ clknet_3_1__leaf_clk reg32_work.bit21.BitData _0058_ VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__dfrtp_2
X_1178_ _0563_ _0564_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__and2b_1
X_1247_ _0148_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1032_ net65 VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__buf_2
X_1101_ _0491_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__buf_2
XFILLER_0_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput40 B[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_0747_ _0268_ _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput62 B[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
Xinput51 B[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
X_0816_ _0330_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_4
X_0678_ _0201_ VGND VGND VPWR VPWR cycle_reg.bit4.BitData sky130_fd_sc_hd__clkbuf_1
X_0601_ _0158_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1015_ _0476_ VGND VGND VPWR VPWR reg32_result.bit29.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ clknet_3_1__leaf_clk _0118_ _0022_ VGND VGND VPWR VPWR reg32_denom.bit16.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_0995_ _0466_ VGND VGND VPWR VPWR reg32_result.bit19.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0780_ _0298_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1194_ _0575_ _0576_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__and2b_1
Xinput5 A[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_1332_ clknet_3_3__leaf_clk reg32_result.bit4.BitData _0074_ VGND VGND VPWR VPWR
+ net93 sky130_fd_sc_hd__dfrtp_1
X_1263_ clknet_3_4__leaf_clk cycle_reg.bit4.BitData _0005_ VGND VGND VPWR VPWR cycle_reg.bit4.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ _0457_ VGND VGND VPWR VPWR reg32_result.bit11.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0832_ _0237_ _0240_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__nor2_1
X_0763_ _0253_ _0262_ _0274_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o31a_2
X_0901_ net162 _0394_ _0404_ _0391_ VGND VGND VPWR VPWR reg32_work.bit19.BitData sky130_fd_sc_hd__o211a_1
X_1315_ clknet_3_0__leaf_clk reg32_work.bit20.BitData _0057_ VGND VGND VPWR VPWR net111
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0694_ reg32_denom.bit18.BitOut net107 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__xnor2_1
X_1177_ _0569_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_1246_ _0140_ _0141_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _0489_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__buf_2
X_1031_ _0190_ _0199_ VGND VGND VPWR VPWR u1.d sky130_fd_sc_hd__nand2_1
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput52 B[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
X_0746_ net128 reg32_denom.bit8.BitOut VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and2b_1
Xinput30 A[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
Xinput41 B[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
X_0815_ _0336_ VGND VGND VPWR VPWR reg32_work.bit1.BitData sky130_fd_sc_hd__clkbuf_1
Xinput63 B[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
X_0677_ _0199_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or2_1
X_1229_ _0138_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0600_ net53 reg32_denom.bit28.BitOut _0154_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1014_ net22 net140 _0191_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
X_0729_ _0249_ net127 _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0994_ net11 net76 _0459_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1331_ clknet_3_2__leaf_clk reg32_result.bit3.BitData _0073_ VGND VGND VPWR VPWR
+ net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 A[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_1193_ _0578_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_1262_ clknet_3_4__leaf_clk cycle_reg.bit3.BitData _0004_ VGND VGND VPWR VPWR cycle_reg.bit3.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ net3 net68 _0448_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0900_ _0347_ _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__nand2_1
X_0831_ _0245_ _0247_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nand2_1
X_0762_ _0262_ _0278_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__o21a_1
X_0693_ reg32_denom.bit19.BitOut net108 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__xor2_1
X_1314_ clknet_3_0__leaf_clk reg32_work.bit19.BitData _0056_ VGND VGND VPWR VPWR net109
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1176_ _0563_ _0564_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and2b_1
X_1245_ _0147_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _0483_ _0488_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__nor2_1
XFILLER_0_33_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 A[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_0814_ _0192_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__and2_1
Xinput31 A[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput64 B[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
Xinput42 B[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
X_0745_ reg32_denom.bit8.BitOut net128 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__and2b_1
Xinput53 B[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
X_0676_ cycle_reg.bit4.BitOut _0197_ net132 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a21o_1
X_1228_ _0587_ _0588_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1159_ _0559_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1013_ _0475_ VGND VGND VPWR VPWR reg32_result.bit28.BitData sky130_fd_sc_hd__clkbuf_1
X_0728_ _0249_ net127 _0241_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o21a_1
X_0659_ net33 reg32_denom.bit0.BitOut _0182_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0465_ VGND VGND VPWR VPWR reg32_result.bit18.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1330_ clknet_3_2__leaf_clk reg32_result.bit2.BitData _0072_ VGND VGND VPWR VPWR
+ net89 sky130_fd_sc_hd__dfrtp_1
X_1261_ clknet_3_4__leaf_clk cycle_reg.bit2.BitData _0003_ VGND VGND VPWR VPWR cycle_reg.bit2.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1192_ _0575_ _0576_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__and2b_1
Xinput7 A[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_0976_ _0456_ VGND VGND VPWR VPWR reg32_result.bit10.BitData sky130_fd_sc_hd__clkbuf_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ net139 _0337_ _0348_ _0190_ VGND VGND VPWR VPWR reg32_work.bit4.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0692_ _0204_ _0207_ _0211_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or4_1
X_0761_ reg32_denom.bit15.BitOut _0279_ _0280_ reg32_denom.bit14.BitOut _0283_ VGND
+ VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1313_ clknet_3_0__leaf_clk reg32_work.bit18.BitData _0055_ VGND VGND VPWR VPWR net108
+ sky130_fd_sc_hd__dfrtp_2
X_1244_ _0140_ _0141_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and2b_1
X_1175_ _0568_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0959_ _0447_ VGND VGND VPWR VPWR reg32_result.bit2.BitData sky130_fd_sc_hd__clkbuf_1
Xoutput130 net130 VGND VGND VPWR VPWR R[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 A[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 A[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput54 B[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XFILLER_0_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput21 A[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput43 B[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
X_0813_ net99 _0334_ net133 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
Xinput65 reset VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
X_0744_ _0263_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__or2_1
X_0675_ net135 _0197_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__nor2_1
X_1227_ _0137_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_1158_ _0551_ _0552_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__and2b_1
X_1089_ _0521_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ net21 net86 _0191_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0727_ _0237_ _0246_ _0245_ _0244_ _0243_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0658_ _0188_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0992_ net10 net75 _0459_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 A[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ _0577_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_1260_ clknet_3_4__leaf_clk cycle_reg.bit1.BitData _0002_ VGND VGND VPWR VPWR cycle_reg.bit1.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ net2 net98 _0448_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ _0281_ _0259_ _0282_ _0256_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o211ai_1
X_0691_ _0212_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1174_ _0563_ _0564_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__and2b_1
X_1312_ clknet_3_1__leaf_clk reg32_work.bit17.BitData _0054_ VGND VGND VPWR VPWR net107
+ sky130_fd_sc_hd__dfrtp_1
X_1243_ _0146_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0958_ net23 net165 _0182_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux2_1
X_0889_ _0221_ _0286_ _0219_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o21ai_1
Xoutput120 net120 VGND VGND VPWR VPWR R[29] sky130_fd_sc_hd__buf_2
Xoutput131 net131 VGND VGND VPWR VPWR err sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput33 B[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput11 A[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_0743_ _0264_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 A[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput55 B[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
Xinput66 start VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xinput44 B[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
X_0812_ _0230_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__xnor2_1
X_0674_ _0197_ _0198_ VGND VGND VPWR VPWR cycle_reg.bit3.BitData sky130_fd_sc_hd__nand2_1
X_1226_ _0587_ _0588_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and2b_1
X_1157_ _0558_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
X_1088_ _0515_ _0516_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1011_ _0474_ VGND VGND VPWR VPWR reg32_result.bit27.BitData sky130_fd_sc_hd__clkbuf_1
X_0726_ reg32_denom.bit7.BitOut VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0657_ net43 reg32_denom.bit19.BitOut _0182_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1209_ _0586_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0709_ reg32_denom.bit1.BitOut net99 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0991_ _0464_ VGND VGND VPWR VPWR reg32_result.bit17.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 A[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_0_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0974_ _0455_ VGND VGND VPWR VPWR reg32_result.bit9.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0690_ reg32_denom.bit22.BitOut net112 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2b_1
X_1311_ clknet_3_1__leaf_clk reg32_work.bit16.BitData _0053_ VGND VGND VPWR VPWR net106
+ sky130_fd_sc_hd__dfrtp_1
X_1173_ _0567_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_1242_ _0140_ _0141_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2b_1
Xoutput121 net121 VGND VGND VPWR VPWR R[2] sky130_fd_sc_hd__clkbuf_4
Xoutput110 net110 VGND VGND VPWR VPWR R[1] sky130_fd_sc_hd__clkbuf_4
Xoutput132 net132 VGND VGND VPWR VPWR ok sky130_fd_sc_hd__clkbuf_4
X_0957_ _0446_ VGND VGND VPWR VPWR reg32_result.bit1.BitData sky130_fd_sc_hd__clkbuf_1
X_0888_ _0330_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput34 B[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
X_0742_ net130 reg32_denom.bit10.BitOut VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__and2b_1
Xinput56 B[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_1
Xinput45 B[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput23 A[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 A[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_0673_ net134 _0195_ net132 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a21oi_1
X_0811_ _0232_ _0231_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or2b_1
X_1225_ _0136_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_1156_ _0551_ _0552_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__and2b_1
X_1087_ _0520_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1010_ net20 net85 _0191_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_0725_ _0243_ _0244_ _0245_ _0247_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0656_ _0187_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1208_ _0575_ _0576_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1139_ _0548_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 cycle_reg.bit3.BitOut VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0639_ _0178_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_0708_ net99 reg32_denom.bit1.BitOut VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0990_ net9 net74 _0459_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ net32 net97 _0448_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ clknet_3_3__leaf_clk reg32_work.bit15.BitData _0052_ VGND VGND VPWR VPWR net105
+ sky130_fd_sc_hd__dfrtp_2
X_1241_ _0145_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_1172_ _0563_ _0564_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ net12 net67 _0182_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
Xoutput111 net111 VGND VGND VPWR VPWR R[20] sky130_fd_sc_hd__clkbuf_4
Xoutput100 net100 VGND VGND VPWR VPWR R[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput122 net122 VGND VGND VPWR VPWR R[30] sky130_fd_sc_hd__clkbuf_4
X_0887_ net153 _0337_ _0393_ _0391_ VGND VGND VPWR VPWR reg32_work.bit16.BitData sky130_fd_sc_hd__o211a_1
Xinput13 A[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_0810_ net157 _0332_ VGND VGND VPWR VPWR reg32_work.bit0.BitData sky130_fd_sc_hd__nor2_1
Xinput24 A[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
X_0741_ reg32_denom.bit10.BitOut net130 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__and2b_1
Xinput46 B[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 B[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
X_0672_ net134 _0195_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__or2_1
Xinput35 B[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
X_1224_ _0587_ _0588_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__and2b_1
X_1155_ _0557_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
X_1086_ _0515_ _0516_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__and2b_1
X_0939_ _0313_ _0317_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0724_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0655_ net54 reg32_denom.bit29.BitOut _0182_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
X_1207_ _0585_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1138_ _0539_ _0540_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1069_ _0510_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 cycle_reg.bit4.BitOut VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0707_ net91 reg32_denom.bit0.BitOut VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__or2b_1
X_0638_ net34 reg32_denom.bit10.BitOut _0171_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0972_ _0454_ VGND VGND VPWR VPWR reg32_result.bit8.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1171_ _0566_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_1240_ _0140_ _0141_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ _0338_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nand2_1
X_0955_ _0445_ VGND VGND VPWR VPWR reg32_result.bit0.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput112 net112 VGND VGND VPWR VPWR R[21] sky130_fd_sc_hd__clkbuf_4
Xoutput123 net123 VGND VGND VPWR VPWR R[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput101 net101 VGND VGND VPWR VPWR R[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 A[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_0740_ reg32_denom.bit11.BitOut net100 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__xor2_1
Xinput25 A[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
Xinput36 B[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput58 B[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
Xinput47 B[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
X_0671_ _0196_ VGND VGND VPWR VPWR cycle_reg.bit2.BitData sky130_fd_sc_hd__clkbuf_1
X_1223_ _0135_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1154_ _0551_ _0552_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2b_1
X_1085_ _0519_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0869_ net101 _0337_ _0379_ _0190_ VGND VGND VPWR VPWR reg32_work.bit12.BitData sky130_fd_sc_hd__o211a_1
X_0938_ _0394_ _0432_ _0433_ VGND VGND VPWR VPWR reg32_work.bit27.BitData sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0723_ reg32_denom.bit5.BitOut net125 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0654_ _0186_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_1137_ _0547_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_1206_ _0575_ _0576_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__and2b_1
X_1068_ _0503_ _0504_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 cycle_reg.bit0.BitOut VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap133 _0329_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_4
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0706_ _0227_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__nand2_1
X_0637_ _0177_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0971_ net31 net96 _0448_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ _0563_ _0564_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__and2b_1
X_0885_ _0221_ _0286_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__xnor2_1
X_0954_ net1 _0330_ _0182_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
Xoutput102 net102 VGND VGND VPWR VPWR R[12] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR R[22] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 VGND VGND VPWR VPWR R[3] sky130_fd_sc_hd__clkbuf_4
X_1299_ clknet_3_4__leaf_clk reg32_work.bit4.BitData _0041_ VGND VGND VPWR VPWR net125
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 B[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput15 A[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 A[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput59 B[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
Xinput48 B[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
X_0670_ _0194_ net132 _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__or3b_1
X_1222_ _0587_ _0588_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__and2b_1
X_1153_ _0556_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_1084_ _0515_ _0516_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0868_ _0377_ _0378_ _0347_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o21ai_1
X_0937_ net117 _0330_ _0192_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o21ai_1
X_0799_ reg32_denom.bit31.BitOut net122 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0722_ net125 reg32_denom.bit5.BitOut VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0653_ net57 reg32_denom.bit31.BitOut _0182_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
X_1136_ _0539_ _0540_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__and2b_1
X_1067_ _0509_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1205_ _0584_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 cycle_reg.bit1.BitOut VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0705_ net110 reg32_denom.bit2.BitOut VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or2b_1
X_0636_ net35 reg32_denom.bit11.BitOut _0171_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1119_ _0537_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0619_ net55 reg32_denom.bit2.BitOut _0160_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
X_0970_ _0453_ VGND VGND VPWR VPWR reg32_result.bit7.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput125 net125 VGND VGND VPWR VPWR R[4] sky130_fd_sc_hd__clkbuf_4
Xoutput103 net103 VGND VGND VPWR VPWR R[13] sky130_fd_sc_hd__clkbuf_4
Xoutput114 net114 VGND VGND VPWR VPWR R[23] sky130_fd_sc_hd__clkbuf_4
X_0953_ _0322_ _0443_ _0444_ VGND VGND VPWR VPWR reg32_work.bit31.BitData sky130_fd_sc_hd__o21a_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0884_ net104 _0337_ _0390_ _0391_ VGND VGND VPWR VPWR reg32_work.bit15.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_37_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1298_ clknet_3_5__leaf_clk reg32_work.bit3.BitData _0040_ VGND VGND VPWR VPWR net124
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput38 B[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
Xinput27 A[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
Xinput49 B[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
Xinput16 A[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_1221_ _0134_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_1152_ _0551_ _0552_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and2b_1
X_1083_ _0518_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
X_0936_ _0298_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0867_ _0278_ _0376_ _0261_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0798_ _0319_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or2_1
X_0721_ reg32_denom.bit7.BitOut net127 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__xnor2_2
X_0652_ _0185_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1204_ _0575_ _0576_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1135_ _0546_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1066_ _0503_ _0504_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and2b_1
X_0919_ _0347_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nand2_1
Xhold5 net118 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0635_ _0176_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0704_ reg32_denom.bit2.BitOut net110 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1118_ _0527_ _0528_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and2b_1
X_1049_ _0499_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0618_ _0167_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0952_ reg32_denom.bit31.BitOut _0319_ _0441_ net122 _0154_ VGND VGND VPWR VPWR _0444_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput104 net104 VGND VGND VPWR VPWR R[14] sky130_fd_sc_hd__buf_2
XFILLER_0_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput126 net126 VGND VGND VPWR VPWR R[5] sky130_fd_sc_hd__buf_2
Xoutput115 net115 VGND VGND VPWR VPWR R[24] sky130_fd_sc_hd__clkbuf_4
X_0883_ _0154_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1297_ clknet_3_4__leaf_clk reg32_work.bit2.BitData _0039_ VGND VGND VPWR VPWR net121
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 A[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
Xinput39 B[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
Xinput17 A[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1220_ _0587_ _0588_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__and2b_1
X_1151_ _0555_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1082_ _0515_ _0516_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and2b_1
X_0866_ _0261_ _0278_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__and3_1
X_0935_ _0302_ _0427_ _0299_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0797_ net120 reg32_denom.bit30.BitOut VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1349_ clknet_3_6__leaf_clk reg32_result.bit21.BitData _0091_ VGND VGND VPWR VPWR
+ net80 sky130_fd_sc_hd__dfrtp_2
X_0720_ _0241_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0651_ net59 reg32_denom.bit4.BitOut _0182_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux2_1
X_1134_ _0539_ _0540_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__and2b_1
X_1203_ _0583_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1065_ _0508_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_0849_ net141 _0337_ _0363_ _0190_ VGND VGND VPWR VPWR reg32_work.bit8.BitData sky130_fd_sc_hd__o211a_1
X_0918_ _0213_ _0416_ _0210_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 net124 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0703_ net121 reg32_denom.bit3.BitOut VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__and2b_1
X_0634_ net36 reg32_denom.bit12.BitOut _0171_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
X_1117_ _0536_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1048_ _0490_ _0492_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0617_ net45 net166 _0160_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0951_ _0319_ _0441_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nor2_1
X_0882_ _0338_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nand2_1
Xoutput116 net116 VGND VGND VPWR VPWR R[25] sky130_fd_sc_hd__clkbuf_4
Xoutput105 net105 VGND VGND VPWR VPWR R[15] sky130_fd_sc_hd__clkbuf_4
Xoutput127 net127 VGND VGND VPWR VPWR R[6] sky130_fd_sc_hd__clkbuf_4
X_1296_ clknet_3_6__leaf_clk reg32_work.bit1.BitData _0038_ VGND VGND VPWR VPWR net110
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 A[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
Xinput29 A[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
X_1150_ _0551_ _0552_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and2b_1
X_1081_ _0517_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
X_0865_ _0253_ _0274_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or2_1
X_0934_ _0430_ VGND VGND VPWR VPWR reg32_work.bit26.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0796_ reg32_denom.bit30.BitOut net120 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__and2b_1
X_1348_ clknet_3_6__leaf_clk reg32_result.bit20.BitData _0090_ VGND VGND VPWR VPWR
+ net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1279_ clknet_3_4__leaf_clk _0117_ _0021_ VGND VGND VPWR VPWR reg32_denom.bit15.BitOut
+ sky130_fd_sc_hd__dfrtp_2
X_0650_ _0184_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_1133_ _0545_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_1064_ _0503_ _0504_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__and2b_1
X_1202_ _0575_ _0576_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0848_ _0338_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__nand2_1
X_0779_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__inv_2
X_0917_ _0213_ _0210_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__and3_1
Xhold7 net87 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0633_ _0175_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_0702_ _0218_ _0221_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1047_ _0498_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_1
X_1116_ _0527_ _0528_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0616_ _0166_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0950_ net145 _0394_ _0442_ _0391_ VGND VGND VPWR VPWR reg32_work.bit30.BitData sky130_fd_sc_hd__o211a_1
X_0881_ _0255_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__xnor2_1
Xoutput128 net128 VGND VGND VPWR VPWR R[7] sky130_fd_sc_hd__clkbuf_4
Xoutput117 net117 VGND VGND VPWR VPWR R[26] sky130_fd_sc_hd__clkbuf_4
Xoutput106 net106 VGND VGND VPWR VPWR R[16] sky130_fd_sc_hd__clkbuf_4
X_1295_ clknet_3_6__leaf_clk net158 _0037_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 A[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_1080_ _0515_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and2b_1
X_0864_ _0375_ VGND VGND VPWR VPWR reg32_work.bit11.BitData sky130_fd_sc_hd__clkbuf_1
X_0933_ _0154_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__and2_1
X_0795_ _0313_ _0316_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nand3_2
XFILLER_0_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1347_ clknet_3_5__leaf_clk reg32_result.bit19.BitData _0089_ VGND VGND VPWR VPWR
+ net77 sky130_fd_sc_hd__dfrtp_4
X_1278_ clknet_3_4__leaf_clk _0116_ _0020_ VGND VGND VPWR VPWR reg32_denom.bit14.BitOut
+ sky130_fd_sc_hd__dfrtp_2
X_1201_ _0582_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1132_ _0539_ _0540_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2b_1
X_1063_ _0507_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_0916_ _0205_ _0203_ _0406_ _0214_ _0202_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a311o_1
X_0847_ _0360_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or2b_1
X_0778_ _0299_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold8 net128 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
X_0632_ net37 reg32_denom.bit13.BitOut _0171_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
X_0701_ _0222_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1115_ _0535_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_1046_ _0490_ _0492_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0615_ net46 reg32_denom.bit21.BitOut _0160_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1029_ _0484_ _0485_ _0486_ _0487_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR R[17] sky130_fd_sc_hd__clkbuf_4
X_0880_ _0254_ _0383_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput129 net129 VGND VGND VPWR VPWR R[8] sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 VGND VGND VPWR VPWR R[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1294_ clknet_3_1__leaf_clk _0132_ _0036_ VGND VGND VPWR VPWR reg32_denom.bit30.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ net116 _0428_ net133 VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ _0192_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and2_1
X_0794_ reg32_denom.bit28.BitOut net118 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__xnor2_2
X_1346_ clknet_3_7__leaf_clk reg32_result.bit18.BitData _0088_ VGND VGND VPWR VPWR
+ net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1277_ clknet_3_4__leaf_clk _0115_ _0019_ VGND VGND VPWR VPWR reg32_denom.bit13.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1200_ _0575_ _0576_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1131_ _0544_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
X_1062_ _0503_ _0504_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0915_ _0415_ VGND VGND VPWR VPWR reg32_work.bit22.BitData sky130_fd_sc_hd__clkbuf_1
X_0846_ _0253_ _0270_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__nand2_1
X_0777_ net116 reg32_denom.bit26.BitOut VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__and2b_1
X_1329_ clknet_3_2__leaf_clk reg32_result.bit1.BitData _0071_ VGND VGND VPWR VPWR
+ net78 sky130_fd_sc_hd__dfrtp_1
Xhold9 net111 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ reg32_denom.bit17.BitOut net106 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0631_ _0174_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_1114_ _0527_ _0528_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1045_ _0497_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0829_ _0240_ _0346_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0614_ _0165_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
X_1028_ net55 net42 net41 net40 VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net119 VGND VGND VPWR VPWR R[28] sky130_fd_sc_hd__clkbuf_4
Xoutput108 net108 VGND VGND VPWR VPWR R[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput90 net90 VGND VGND VPWR VPWR D[30] sky130_fd_sc_hd__clkbuf_4
X_1293_ clknet_3_1__leaf_clk _0131_ _0035_ VGND VGND VPWR VPWR reg32_denom.bit3.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ net100 _0373_ net133 VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_1
X_0931_ _0301_ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__xnor2_1
X_0793_ _0314_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__and2b_1
X_1345_ clknet_3_7__leaf_clk reg32_result.bit17.BitData _0087_ VGND VGND VPWR VPWR
+ net75 sky130_fd_sc_hd__dfrtp_1
X_1276_ clknet_3_6__leaf_clk _0114_ _0018_ VGND VGND VPWR VPWR reg32_denom.bit12.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1130_ _0539_ _0540_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1061_ _0506_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
X_0845_ _0253_ _0270_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
X_0914_ _0154_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and2_1
X_0776_ reg32_denom.bit26.BitOut net116 VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1328_ clknet_3_3__leaf_clk reg32_result.bit0.BitData _0070_ VGND VGND VPWR VPWR
+ net67 sky130_fd_sc_hd__dfrtp_2
X_1259_ clknet_3_4__leaf_clk cycle_reg.bit0.BitData _0001_ VGND VGND VPWR VPWR cycle_reg.bit0.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0630_ net38 reg32_denom.bit14.BitOut _0171_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ _0534_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
X_1044_ _0490_ _0492_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0828_ net133 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0759_ _0254_ _0255_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0613_ net47 reg32_denom.bit22.BitOut _0160_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1027_ net48 net47 net46 net45 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR R[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput80 net80 VGND VGND VPWR VPWR D[21] sky130_fd_sc_hd__clkbuf_4
Xoutput91 net91 VGND VGND VPWR VPWR D[31] sky130_fd_sc_hd__clkbuf_4
X_1292_ clknet_3_1__leaf_clk _0130_ _0034_ VGND VGND VPWR VPWR reg32_denom.bit28.BitOut
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0861_ _0263_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__xnor2_1
X_0930_ _0307_ _0308_ _0420_ _0311_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a31o_1
X_0792_ reg32_denom.bit29.BitOut net119 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or2b_1
X_1344_ clknet_3_7__leaf_clk reg32_result.bit16.BitData _0086_ VGND VGND VPWR VPWR
+ net74 sky130_fd_sc_hd__dfrtp_1
X_1275_ clknet_3_6__leaf_clk _0113_ _0017_ VGND VGND VPWR VPWR reg32_denom.bit11.BitOut
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1060_ _0503_ _0504_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0844_ net127 _0337_ _0359_ _0190_ VGND VGND VPWR VPWR reg32_work.bit7.BitData sky130_fd_sc_hd__o211a_1
X_0775_ _0296_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and2b_1
X_0913_ net112 _0413_ _0329_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_1327_ clknet_3_1__leaf_clk _0133_ _0069_ VGND VGND VPWR VPWR reg32_denom.bit9.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_1189_ _0491_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__buf_2
X_1258_ clknet_3_4__leaf_clk u1.d _0000_ VGND VGND VPWR VPWR u1.q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1112_ _0527_ _0528_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__and2b_1
X_1043_ _0496_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ _0236_ _0239_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0758_ _0257_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__inv_2
X_0689_ net112 reg32_denom.bit22.BitOut VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0612_ _0164_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1026_ net64 net56 net58 net53 VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ _0473_ VGND VGND VPWR VPWR reg32_result.bit26.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput70 net70 VGND VGND VPWR VPWR D[12] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR D[3] sky130_fd_sc_hd__clkbuf_4
Xoutput81 net81 VGND VGND VPWR VPWR D[22] sky130_fd_sc_hd__buf_2
X_1291_ clknet_3_2__leaf_clk _0129_ _0033_ VGND VGND VPWR VPWR reg32_denom.bit27.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0860_ _0371_ _0367_ _0264_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21o_1
X_0791_ net119 reg32_denom.bit29.BitOut VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1343_ clknet_3_5__leaf_clk reg32_result.bit15.BitData _0085_ VGND VGND VPWR VPWR
+ net73 sky130_fd_sc_hd__dfrtp_1
X_1274_ clknet_3_6__leaf_clk _0112_ _0016_ VGND VGND VPWR VPWR reg32_denom.bit10.BitOut
+ sky130_fd_sc_hd__dfrtp_1
X_0989_ _0463_ VGND VGND VPWR VPWR reg32_result.bit16.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0912_ _0214_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__xor2_1
X_0843_ _0338_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__nand2_1
X_0774_ net117 reg32_denom.bit27.BitOut VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ clknet_3_0__leaf_clk reg32_work.bit31.BitData _0068_ VGND VGND VPWR VPWR net123
+ sky130_fd_sc_hd__dfrtp_1
X_1188_ _0489_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_2
X_1257_ _0153_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1111_ _0533_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
X_1042_ _0490_ _0492_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0826_ net150 _0337_ _0345_ _0190_ VGND VGND VPWR VPWR reg32_work.bit3.BitData sky130_fd_sc_hd__o211a_1
X_0757_ reg32_denom.bit15.BitOut _0279_ net103 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0688_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1309_ clknet_3_3__leaf_clk reg32_work.bit14.BitData _0051_ VGND VGND VPWR VPWR net104
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0611_ net48 reg32_denom.bit23.BitOut _0160_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
X_1025_ net52 net51 net50 net49 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0809_ reg32_denom.bit0.BitOut net91 _0330_ net132 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ net19 net151 _0191_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput71 net71 VGND VGND VPWR VPWR D[13] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 VGND VGND VPWR VPWR D[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput93 net93 VGND VGND VPWR VPWR D[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1290_ clknet_3_2__leaf_clk _0128_ _0032_ VGND VGND VPWR VPWR reg32_denom.bit26.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ _0295_ _0309_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1342_ clknet_3_5__leaf_clk reg32_result.bit14.BitData _0084_ VGND VGND VPWR VPWR
+ net72 sky130_fd_sc_hd__dfrtp_1
X_1273_ clknet_3_6__leaf_clk _0111_ _0015_ VGND VGND VPWR VPWR reg32_denom.bit1.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0988_ net8 net73 _0459_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0842_ _0244_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__xnor2_1
X_0911_ _0205_ _0203_ _0406_ _0202_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a31o_1
X_0773_ reg32_denom.bit27.BitOut net117 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__and2b_1
X_1325_ clknet_3_0__leaf_clk reg32_work.bit30.BitData _0067_ VGND VGND VPWR VPWR net122
+ sky130_fd_sc_hd__dfrtp_2
X_1256_ _0489_ _0491_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__and2b_1
X_1187_ _0574_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1110_ _0527_ _0528_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1041_ _0495_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0825_ _0338_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0687_ _0208_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0756_ net104 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1239_ _0144_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_1308_ clknet_3_6__leaf_clk reg32_work.bit13.BitData _0050_ VGND VGND VPWR VPWR net103
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0610_ _0163_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
X_1024_ _0479_ _0480_ _0481_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0808_ net156 _0330_ net91 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a21oi_1
X_0739_ _0254_ _0255_ _0258_ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _0472_ VGND VGND VPWR VPWR reg32_result.bit25.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput72 net72 VGND VGND VPWR VPWR D[14] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR D[5] sky130_fd_sc_hd__clkbuf_4
Xoutput83 net83 VGND VGND VPWR VPWR D[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1341_ clknet_3_5__leaf_clk reg32_result.bit13.BitData _0083_ VGND VGND VPWR VPWR
+ net71 sky130_fd_sc_hd__dfrtp_1
X_1272_ clknet_3_6__leaf_clk _0110_ _0014_ VGND VGND VPWR VPWR reg32_denom.bit8.BitOut
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0987_ _0462_ VGND VGND VPWR VPWR reg32_result.bit15.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0841_ _0243_ _0353_ _0241_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a21o_1
X_0772_ _0215_ _0225_ _0286_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o31ai_2
X_0910_ net142 _0394_ _0411_ _0391_ VGND VGND VPWR VPWR reg32_work.bit21.BitData sky130_fd_sc_hd__o211a_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1324_ clknet_3_3__leaf_clk reg32_work.bit29.BitData _0066_ VGND VGND VPWR VPWR net120
+ sky130_fd_sc_hd__dfrtp_2
X_1186_ _0563_ _0564_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__and2b_1
X_1255_ _0152_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1040_ _0490_ _0492_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__and2b_1
X_0755_ reg32_denom.bit11.BitOut _0275_ _0267_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0824_ _0341_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__xnor2_1
X_0686_ reg32_denom.bit23.BitOut net113 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2b_1
X_1307_ clknet_3_7__leaf_clk reg32_work.bit12.BitData _0049_ VGND VGND VPWR VPWR net102
+ sky130_fd_sc_hd__dfrtp_2
X_1169_ _0565_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_1238_ _0140_ _0141_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1023_ net57 net54 net43 net33 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or4_1
X_0807_ net133 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_4
X_0738_ _0259_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__or2_1
X_0669_ cycle_reg.bit0.BitOut cycle_reg.bit1.BitOut cycle_reg.bit2.BitOut VGND VGND
+ VPWR VPWR _0195_ sky130_fd_sc_hd__or3_1
XANTENNA_3 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ net18 net83 _0191_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput73 net73 VGND VGND VPWR VPWR D[15] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 VGND VGND VPWR VPWR D[6] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR D[25] sky130_fd_sc_hd__buf_2
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1340_ clknet_3_7__leaf_clk reg32_result.bit12.BitData _0082_ VGND VGND VPWR VPWR
+ net70 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1271_ clknet_3_4__leaf_clk _0109_ _0013_ VGND VGND VPWR VPWR reg32_denom.bit7.BitOut
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0986_ net7 net147 _0459_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0840_ _0356_ VGND VGND VPWR VPWR reg32_work.bit6.BitData sky130_fd_sc_hd__clkbuf_1
X_0771_ _0293_ _0213_ _0209_ _0208_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a31o_1
X_1323_ clknet_3_3__leaf_clk reg32_work.bit28.BitData _0065_ VGND VGND VPWR VPWR net119
+ sky130_fd_sc_hd__dfrtp_2
X_1185_ _0573_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_1254_ _0489_ _0491_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0969_ net30 net95 _0448_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0754_ reg32_denom.bit11.BitOut _0275_ _0264_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a21bo_1
X_0685_ net113 reg32_denom.bit23.BitOut VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0823_ _0342_ _0226_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__nor2_1
X_1306_ clknet_3_7__leaf_clk reg32_work.bit11.BitData _0048_ VGND VGND VPWR VPWR net101
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1168_ _0563_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and2b_1
X_1099_ _0526_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
X_1237_ _0143_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1022_ net62 net61 net60 net59 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0806_ _0318_ _0323_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o21ai_2
X_0668_ cycle_reg.bit0.BitOut cycle_reg.bit1.BitOut cycle_reg.bit2.BitOut VGND VGND
+ VPWR VPWR _0194_ sky130_fd_sc_hd__o21a_1
X_0737_ net101 reg32_denom.bit12.BitOut VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_0599_ _0157_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1005_ _0471_ VGND VGND VPWR VPWR reg32_result.bit24.BitData sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput85 net85 VGND VGND VPWR VPWR D[26] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 VGND VGND VPWR VPWR D[7] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR D[16] sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

