magic
tech sky130A
magscale 1 2
timestamp 1700823269
<< viali >>
rect 1593 26537 1627 26571
rect 2237 26537 2271 26571
rect 7389 26537 7423 26571
rect 9137 26537 9171 26571
rect 11069 26537 11103 26571
rect 11897 26537 11931 26571
rect 14473 26537 14507 26571
rect 17049 26537 17083 26571
rect 19441 26537 19475 26571
rect 20269 26537 20303 26571
rect 20913 26537 20947 26571
rect 23949 26537 23983 26571
rect 3801 26469 3835 26503
rect 9965 26469 9999 26503
rect 15577 26469 15611 26503
rect 17509 26469 17543 26503
rect 18337 26469 18371 26503
rect 22569 26469 22603 26503
rect 2697 26401 2731 26435
rect 24593 26401 24627 26435
rect 2973 26333 3007 26367
rect 3985 26333 4019 26367
rect 5273 26333 5307 26367
rect 5917 26333 5951 26367
rect 6561 26333 6595 26367
rect 9505 26333 9539 26367
rect 9781 26333 9815 26367
rect 12357 26333 12391 26367
rect 13001 26333 13035 26367
rect 15761 26333 15795 26367
rect 16957 26333 16991 26367
rect 17693 26333 17727 26367
rect 18153 26333 18187 26367
rect 22385 26333 22419 26367
rect 23213 26333 23247 26367
rect 23305 26333 23339 26367
rect 24869 26333 24903 26367
rect 1501 26265 1535 26299
rect 2145 26265 2179 26299
rect 7297 26265 7331 26299
rect 9045 26265 9079 26299
rect 10977 26265 11011 26299
rect 11805 26265 11839 26299
rect 14381 26265 14415 26299
rect 15025 26265 15059 26299
rect 19349 26265 19383 26299
rect 20177 26265 20211 26299
rect 20821 26265 20855 26299
rect 21925 26265 21959 26299
rect 23857 26265 23891 26299
rect 5457 26197 5491 26231
rect 6101 26197 6135 26231
rect 6745 26197 6779 26231
rect 9689 26197 9723 26231
rect 12541 26197 12575 26231
rect 13185 26197 13219 26231
rect 15117 26197 15151 26231
rect 22017 26197 22051 26231
rect 23029 26197 23063 26231
rect 23489 26197 23523 26231
rect 1961 25993 1995 26027
rect 7849 25993 7883 26027
rect 7941 25993 7975 26027
rect 16313 25993 16347 26027
rect 17601 25993 17635 26027
rect 21005 25993 21039 26027
rect 18153 25925 18187 25959
rect 24225 25925 24259 25959
rect 1869 25857 1903 25891
rect 2421 25857 2455 25891
rect 2881 25857 2915 25891
rect 3157 25857 3191 25891
rect 10241 25857 10275 25891
rect 11713 25857 11747 25891
rect 11989 25857 12023 25891
rect 16221 25857 16255 25891
rect 16405 25857 16439 25891
rect 17785 25857 17819 25891
rect 21649 25857 21683 25891
rect 23765 25857 23799 25891
rect 24593 25857 24627 25891
rect 8125 25789 8159 25823
rect 8309 25789 8343 25823
rect 8585 25789 8619 25823
rect 10057 25789 10091 25823
rect 10885 25789 10919 25823
rect 17877 25789 17911 25823
rect 19625 25789 19659 25823
rect 21097 25789 21131 25823
rect 21189 25789 21223 25823
rect 24685 25789 24719 25823
rect 24961 25789 24995 25823
rect 11253 25721 11287 25755
rect 2513 25653 2547 25687
rect 3065 25653 3099 25687
rect 3341 25653 3375 25687
rect 7481 25653 7515 25687
rect 10793 25653 10827 25687
rect 11345 25653 11379 25687
rect 11529 25653 11563 25687
rect 11805 25653 11839 25687
rect 20637 25653 20671 25687
rect 21465 25653 21499 25687
rect 23949 25653 23983 25687
rect 1593 25449 1627 25483
rect 8217 25449 8251 25483
rect 8953 25449 8987 25483
rect 9781 25449 9815 25483
rect 12541 25449 12575 25483
rect 15853 25449 15887 25483
rect 16865 25449 16899 25483
rect 17417 25449 17451 25483
rect 17877 25449 17911 25483
rect 18797 25449 18831 25483
rect 20361 25449 20395 25483
rect 24869 25449 24903 25483
rect 25421 25449 25455 25483
rect 9597 25381 9631 25415
rect 13001 25381 13035 25415
rect 13185 25381 13219 25415
rect 19625 25381 19659 25415
rect 20177 25381 20211 25415
rect 6469 25313 6503 25347
rect 10425 25313 10459 25347
rect 11069 25313 11103 25347
rect 14105 25313 14139 25347
rect 18521 25313 18555 25347
rect 19717 25313 19751 25347
rect 1961 25245 1995 25279
rect 6377 25245 6411 25279
rect 8493 25245 8527 25279
rect 8769 25245 8803 25279
rect 9137 25245 9171 25279
rect 10793 25245 10827 25279
rect 13921 25245 13955 25279
rect 16129 25245 16163 25279
rect 16773 25245 16807 25279
rect 17325 25245 17359 25279
rect 18245 25245 18279 25279
rect 18981 25245 19015 25279
rect 20453 25245 20487 25279
rect 24225 25245 24259 25279
rect 24685 25245 24719 25279
rect 1501 25177 1535 25211
rect 6745 25177 6779 25211
rect 9229 25177 9263 25211
rect 10241 25177 10275 25211
rect 12725 25177 12759 25211
rect 14381 25177 14415 25211
rect 19257 25177 19291 25211
rect 19901 25177 19935 25211
rect 20729 25177 20763 25211
rect 25145 25177 25179 25211
rect 2145 25109 2179 25143
rect 6193 25109 6227 25143
rect 8309 25109 8343 25143
rect 8585 25109 8619 25143
rect 9689 25109 9723 25143
rect 10149 25109 10183 25143
rect 13737 25109 13771 25143
rect 16681 25109 16715 25143
rect 17233 25109 17267 25143
rect 17785 25109 17819 25143
rect 18337 25109 18371 25143
rect 22201 25109 22235 25143
rect 24041 25109 24075 25143
rect 6377 24905 6411 24939
rect 11989 24905 12023 24939
rect 13185 24905 13219 24939
rect 15117 24905 15151 24939
rect 16405 24905 16439 24939
rect 17141 24905 17175 24939
rect 21465 24905 21499 24939
rect 6745 24837 6779 24871
rect 7665 24837 7699 24871
rect 9137 24837 9171 24871
rect 12725 24837 12759 24871
rect 16681 24837 16715 24871
rect 6837 24769 6871 24803
rect 8217 24769 8251 24803
rect 8861 24769 8895 24803
rect 12449 24769 12483 24803
rect 15393 24769 15427 24803
rect 15485 24769 15519 24803
rect 15577 24769 15611 24803
rect 15761 24769 15795 24803
rect 16037 24769 16071 24803
rect 21373 24769 21407 24803
rect 21649 24769 21683 24803
rect 7021 24701 7055 24735
rect 7757 24701 7791 24735
rect 7941 24701 7975 24735
rect 10885 24701 10919 24735
rect 11529 24701 11563 24735
rect 13277 24701 13311 24735
rect 13553 24701 13587 24735
rect 16129 24701 16163 24735
rect 17233 24701 17267 24735
rect 17693 24701 17727 24735
rect 17785 24701 17819 24735
rect 19349 24701 19383 24735
rect 19625 24701 19659 24735
rect 21097 24701 21131 24735
rect 8769 24633 8803 24667
rect 11897 24633 11931 24667
rect 13001 24633 13035 24667
rect 15025 24633 15059 24667
rect 16957 24633 16991 24667
rect 17601 24633 17635 24667
rect 18153 24633 18187 24667
rect 21189 24633 21223 24667
rect 7297 24565 7331 24599
rect 12265 24565 12299 24599
rect 18245 24565 18279 24599
rect 8125 24361 8159 24395
rect 10425 24361 10459 24395
rect 14105 24361 14139 24395
rect 15301 24361 15335 24395
rect 15945 24361 15979 24395
rect 17509 24361 17543 24395
rect 20177 24361 20211 24395
rect 10241 24293 10275 24327
rect 13093 24293 13127 24327
rect 16497 24293 16531 24327
rect 20085 24293 20119 24327
rect 20637 24293 20671 24327
rect 10333 24225 10367 24259
rect 11345 24225 11379 24259
rect 13369 24225 13403 24259
rect 14933 24225 14967 24259
rect 16589 24225 16623 24259
rect 17601 24225 17635 24259
rect 20821 24225 20855 24259
rect 8309 24157 8343 24191
rect 10609 24157 10643 24191
rect 13921 24157 13955 24191
rect 14381 24157 14415 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15025 24157 15059 24191
rect 15209 24157 15243 24191
rect 15393 24157 15427 24191
rect 15669 24157 15703 24191
rect 16405 24157 16439 24191
rect 16681 24157 16715 24191
rect 16865 24157 16899 24191
rect 17325 24157 17359 24191
rect 17417 24157 17451 24191
rect 19717 24157 19751 24191
rect 20361 24157 20395 24191
rect 21373 24157 21407 24191
rect 21649 24157 21683 24191
rect 25237 24157 25271 24191
rect 1501 24089 1535 24123
rect 9873 24089 9907 24123
rect 11621 24089 11655 24123
rect 17049 24089 17083 24123
rect 1593 24021 1627 24055
rect 16129 24021 16163 24055
rect 16221 24021 16255 24055
rect 17233 24021 17267 24055
rect 21189 24021 21223 24055
rect 21465 24021 21499 24055
rect 25421 24021 25455 24055
rect 9413 23817 9447 23851
rect 12265 23817 12299 23851
rect 13737 23817 13771 23851
rect 15853 23817 15887 23851
rect 16129 23817 16163 23851
rect 17049 23817 17083 23851
rect 20177 23817 20211 23851
rect 20913 23817 20947 23851
rect 11805 23749 11839 23783
rect 22109 23749 22143 23783
rect 1409 23681 1443 23715
rect 5549 23681 5583 23715
rect 6561 23681 6595 23715
rect 8217 23681 8251 23715
rect 8401 23681 8435 23715
rect 9643 23681 9677 23715
rect 9781 23681 9815 23715
rect 9873 23681 9907 23715
rect 10057 23681 10091 23715
rect 10333 23681 10367 23715
rect 13921 23681 13955 23715
rect 15761 23681 15795 23715
rect 15945 23681 15979 23715
rect 16043 23681 16077 23715
rect 16221 23681 16255 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 19809 23681 19843 23715
rect 19993 23681 20027 23715
rect 20361 23681 20395 23715
rect 20729 23681 20763 23715
rect 21281 23681 21315 23715
rect 21833 23681 21867 23715
rect 25329 23681 25363 23715
rect 5825 23613 5859 23647
rect 6469 23613 6503 23647
rect 8309 23613 8343 23647
rect 21373 23613 21407 23647
rect 21557 23613 21591 23647
rect 1593 23545 1627 23579
rect 5365 23545 5399 23579
rect 6929 23545 6963 23579
rect 12173 23545 12207 23579
rect 5733 23477 5767 23511
rect 10149 23477 10183 23511
rect 16865 23477 16899 23511
rect 20545 23477 20579 23511
rect 23581 23477 23615 23511
rect 25513 23477 25547 23511
rect 20361 23273 20395 23307
rect 20913 23273 20947 23307
rect 4537 23205 4571 23239
rect 5181 23205 5215 23239
rect 19533 23205 19567 23239
rect 20177 23205 20211 23239
rect 4813 23137 4847 23171
rect 6377 23137 6411 23171
rect 6653 23137 6687 23171
rect 8953 23137 8987 23171
rect 10977 23137 11011 23171
rect 12817 23137 12851 23171
rect 19257 23137 19291 23171
rect 19901 23137 19935 23171
rect 21465 23137 21499 23171
rect 21833 23137 21867 23171
rect 4261 23069 4295 23103
rect 5552 23069 5586 23103
rect 5641 23069 5675 23103
rect 5825 23069 5859 23103
rect 5917 23069 5951 23103
rect 6285 23069 6319 23103
rect 6745 23069 6779 23103
rect 7021 23069 7055 23103
rect 12357 23069 12391 23103
rect 12541 23069 12575 23103
rect 12633 23069 12667 23103
rect 14289 23069 14323 23103
rect 16681 23069 16715 23103
rect 16957 23069 16991 23103
rect 17049 23069 17083 23103
rect 17509 23069 17543 23103
rect 20545 23069 20579 23103
rect 6929 23001 6963 23035
rect 9229 23001 9263 23035
rect 17233 23001 17267 23035
rect 17601 23001 17635 23035
rect 4721 22933 4755 22967
rect 5273 22933 5307 22967
rect 5365 22933 5399 22967
rect 7113 22933 7147 22967
rect 7297 22933 7331 22967
rect 12173 22933 12207 22967
rect 14105 22933 14139 22967
rect 16497 22933 16531 22967
rect 16865 22933 16899 22967
rect 17417 22933 17451 22967
rect 19717 22933 19751 22967
rect 20729 22933 20763 22967
rect 21281 22933 21315 22967
rect 21373 22933 21407 22967
rect 22385 22933 22419 22967
rect 3341 22729 3375 22763
rect 6101 22729 6135 22763
rect 7573 22729 7607 22763
rect 8401 22729 8435 22763
rect 10241 22729 10275 22763
rect 13737 22729 13771 22763
rect 14197 22729 14231 22763
rect 15025 22729 15059 22763
rect 17785 22729 17819 22763
rect 21465 22729 21499 22763
rect 11897 22661 11931 22695
rect 17877 22661 17911 22695
rect 1501 22593 1535 22627
rect 2605 22593 2639 22627
rect 3433 22593 3467 22627
rect 4445 22593 4479 22627
rect 4721 22593 4755 22627
rect 5089 22593 5123 22627
rect 6009 22593 6043 22627
rect 6653 22593 6687 22627
rect 7481 22593 7515 22627
rect 8033 22593 8067 22627
rect 8125 22593 8159 22627
rect 8309 22593 8343 22627
rect 8585 22593 8619 22627
rect 11621 22593 11655 22627
rect 14105 22593 14139 22627
rect 14841 22593 14875 22627
rect 16129 22593 16163 22627
rect 16865 22593 16899 22627
rect 18061 22593 18095 22627
rect 19625 22593 19659 22627
rect 25513 22593 25547 22627
rect 3525 22525 3559 22559
rect 3801 22525 3835 22559
rect 5365 22525 5399 22559
rect 5825 22525 5859 22559
rect 6745 22525 6779 22559
rect 7665 22525 7699 22559
rect 9781 22525 9815 22559
rect 13645 22525 13679 22559
rect 14289 22525 14323 22559
rect 14657 22525 14691 22559
rect 16221 22525 16255 22559
rect 16773 22525 16807 22559
rect 17233 22525 17267 22559
rect 17325 22525 17359 22559
rect 18245 22525 18279 22559
rect 19717 22525 19751 22559
rect 19993 22525 20027 22559
rect 2973 22457 3007 22491
rect 7021 22457 7055 22491
rect 7113 22457 7147 22491
rect 10149 22457 10183 22491
rect 16497 22457 16531 22491
rect 17693 22457 17727 22491
rect 1593 22389 1627 22423
rect 2421 22389 2455 22423
rect 4537 22389 4571 22423
rect 19441 22389 19475 22423
rect 25329 22389 25363 22423
rect 2132 22185 2166 22219
rect 3617 22185 3651 22219
rect 3801 22185 3835 22219
rect 5457 22185 5491 22219
rect 7113 22185 7147 22219
rect 12357 22185 12391 22219
rect 14362 22185 14396 22219
rect 15945 22185 15979 22219
rect 21097 22185 21131 22219
rect 9045 22117 9079 22151
rect 12081 22117 12115 22151
rect 13001 22117 13035 22151
rect 13553 22117 13587 22151
rect 4353 22049 4387 22083
rect 6469 22049 6503 22083
rect 9229 22049 9263 22083
rect 12265 22049 12299 22083
rect 16497 22049 16531 22083
rect 17049 22049 17083 22083
rect 17693 22049 17727 22083
rect 18981 22049 19015 22083
rect 19257 22049 19291 22083
rect 1869 21981 1903 22015
rect 4721 21981 4755 22015
rect 5733 21981 5767 22015
rect 6101 21981 6135 22015
rect 6193 21981 6227 22015
rect 6653 21981 6687 22015
rect 7021 21981 7055 22015
rect 7113 21981 7147 22015
rect 7297 21981 7331 22015
rect 8401 21981 8435 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 8769 21981 8803 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 11345 21981 11379 22015
rect 11805 21981 11839 22015
rect 12541 21981 12575 22015
rect 14105 21981 14139 22015
rect 16313 21981 16347 22015
rect 16773 21981 16807 22015
rect 16957 21981 16991 22015
rect 17141 21981 17175 22015
rect 17325 21981 17359 22015
rect 17785 21981 17819 22015
rect 18705 21981 18739 22015
rect 21281 21981 21315 22015
rect 25513 21981 25547 22015
rect 4169 21913 4203 21947
rect 8125 21913 8159 21947
rect 9505 21913 9539 21947
rect 12725 21913 12759 21947
rect 13277 21913 13311 21947
rect 16405 21913 16439 21947
rect 19533 21913 19567 21947
rect 4261 21845 4295 21879
rect 5273 21845 5307 21879
rect 5825 21845 5859 21879
rect 5917 21845 5951 21879
rect 6929 21845 6963 21879
rect 10977 21845 11011 21879
rect 11161 21845 11195 21879
rect 13185 21845 13219 21879
rect 13737 21845 13771 21879
rect 15853 21845 15887 21879
rect 17509 21845 17543 21879
rect 18153 21845 18187 21879
rect 18337 21845 18371 21879
rect 18797 21845 18831 21879
rect 21005 21845 21039 21879
rect 25329 21845 25363 21879
rect 2145 21641 2179 21675
rect 9137 21641 9171 21675
rect 10517 21641 10551 21675
rect 13277 21641 13311 21675
rect 17325 21641 17359 21675
rect 17877 21641 17911 21675
rect 18613 21641 18647 21675
rect 20085 21641 20119 21675
rect 23857 21641 23891 21675
rect 4721 21573 4755 21607
rect 5733 21573 5767 21607
rect 6377 21573 6411 21607
rect 7113 21573 7147 21607
rect 7389 21573 7423 21607
rect 16681 21573 16715 21607
rect 1501 21505 1535 21539
rect 2329 21505 2363 21539
rect 2421 21505 2455 21539
rect 4629 21505 4663 21539
rect 4813 21505 4847 21539
rect 5917 21505 5951 21539
rect 6101 21505 6135 21539
rect 6193 21505 6227 21539
rect 6561 21505 6595 21539
rect 6837 21505 6871 21539
rect 7021 21505 7055 21539
rect 7297 21505 7331 21539
rect 7481 21505 7515 21539
rect 7849 21505 7883 21539
rect 13461 21505 13495 21539
rect 13553 21505 13587 21539
rect 16313 21505 16347 21539
rect 16405 21505 16439 21539
rect 17141 21505 17175 21539
rect 18797 21505 18831 21539
rect 20453 21505 20487 21539
rect 21649 21505 21683 21539
rect 2697 21437 2731 21471
rect 4169 21437 4203 21471
rect 5181 21437 5215 21471
rect 6653 21437 6687 21471
rect 10057 21437 10091 21471
rect 13829 21437 13863 21471
rect 17049 21437 17083 21471
rect 17417 21437 17451 21471
rect 20545 21437 20579 21471
rect 20637 21437 20671 21471
rect 23949 21437 23983 21471
rect 24133 21437 24167 21471
rect 5549 21369 5583 21403
rect 5641 21369 5675 21403
rect 6745 21369 6779 21403
rect 10333 21369 10367 21403
rect 15301 21369 15335 21403
rect 17693 21369 17727 21403
rect 1593 21301 1627 21335
rect 21465 21301 21499 21335
rect 23489 21301 23523 21335
rect 2697 21097 2731 21131
rect 3341 21097 3375 21131
rect 5457 21097 5491 21131
rect 11253 21097 11287 21131
rect 11621 21097 11655 21131
rect 13645 21097 13679 21131
rect 17141 21097 17175 21131
rect 20821 21097 20855 21131
rect 2605 21029 2639 21063
rect 3157 21029 3191 21063
rect 5641 21029 5675 21063
rect 10057 21029 10091 21063
rect 10517 21029 10551 21063
rect 12173 21029 12207 21063
rect 20637 21029 20671 21063
rect 25513 21029 25547 21063
rect 3249 20961 3283 20995
rect 1409 20893 1443 20927
rect 3525 20893 3559 20927
rect 5181 20893 5215 20927
rect 8769 20893 8803 20927
rect 8953 20893 8987 20927
rect 13829 20893 13863 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 14657 20893 14691 20927
rect 14841 20893 14875 20927
rect 15669 20893 15703 20927
rect 20913 20893 20947 20927
rect 25329 20893 25363 20927
rect 2237 20825 2271 20859
rect 2789 20825 2823 20859
rect 9689 20825 9723 20859
rect 10241 20825 10275 20859
rect 11161 20825 11195 20859
rect 11529 20825 11563 20859
rect 11897 20825 11931 20859
rect 20361 20825 20395 20859
rect 21189 20825 21223 20859
rect 1593 20757 1627 20791
rect 8585 20757 8619 20791
rect 9597 20757 9631 20791
rect 10149 20757 10183 20791
rect 10701 20757 10735 20791
rect 12357 20757 12391 20791
rect 14197 20757 14231 20791
rect 22661 20757 22695 20791
rect 2881 20553 2915 20587
rect 11253 20553 11287 20587
rect 12357 20553 12391 20587
rect 12817 20553 12851 20587
rect 21373 20553 21407 20587
rect 21833 20553 21867 20587
rect 22293 20553 22327 20587
rect 15853 20485 15887 20519
rect 3709 20417 3743 20451
rect 3985 20417 4019 20451
rect 7481 20417 7515 20451
rect 7573 20417 7607 20451
rect 7665 20417 7699 20451
rect 7849 20417 7883 20451
rect 8401 20417 8435 20451
rect 10517 20417 10551 20451
rect 11069 20417 11103 20451
rect 11529 20417 11563 20451
rect 13001 20417 13035 20451
rect 16037 20417 16071 20451
rect 16221 20417 16255 20451
rect 18429 20417 18463 20451
rect 20361 20417 20395 20451
rect 21557 20417 21591 20451
rect 22201 20417 22235 20451
rect 23765 20417 23799 20451
rect 2421 20349 2455 20383
rect 2973 20349 3007 20383
rect 3433 20349 3467 20383
rect 12449 20349 12483 20383
rect 12633 20349 12667 20383
rect 22385 20349 22419 20383
rect 2789 20281 2823 20315
rect 3249 20281 3283 20315
rect 10333 20281 10367 20315
rect 11989 20281 12023 20315
rect 3525 20213 3559 20247
rect 3801 20213 3835 20247
rect 7205 20213 7239 20247
rect 8658 20213 8692 20247
rect 10149 20213 10183 20247
rect 11713 20213 11747 20247
rect 18613 20213 18647 20247
rect 20545 20213 20579 20247
rect 23581 20213 23615 20247
rect 3801 20009 3835 20043
rect 4629 20009 4663 20043
rect 7021 20009 7055 20043
rect 7757 20009 7791 20043
rect 8953 20009 8987 20043
rect 13277 20009 13311 20043
rect 15025 20009 15059 20043
rect 16773 20009 16807 20043
rect 25421 20009 25455 20043
rect 5181 19941 5215 19975
rect 6285 19941 6319 19975
rect 6837 19941 6871 19975
rect 15669 19941 15703 19975
rect 18889 19941 18923 19975
rect 19533 19941 19567 19975
rect 20821 19941 20855 19975
rect 21373 19941 21407 19975
rect 1777 19873 1811 19907
rect 4353 19873 4387 19907
rect 4721 19873 4755 19907
rect 6561 19873 6595 19907
rect 7849 19873 7883 19907
rect 11529 19873 11563 19907
rect 15117 19873 15151 19907
rect 15945 19873 15979 19907
rect 18521 19873 18555 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 21557 19873 21591 19907
rect 24133 19873 24167 19907
rect 4169 19805 4203 19839
rect 4629 19805 4663 19839
rect 4905 19805 4939 19839
rect 5365 19805 5399 19839
rect 6009 19805 6043 19839
rect 7113 19805 7147 19839
rect 7297 19805 7331 19839
rect 7481 19805 7515 19839
rect 7573 19805 7607 19839
rect 7665 19805 7699 19839
rect 8309 19805 8343 19839
rect 8493 19805 8527 19839
rect 9229 19805 9263 19839
rect 9321 19805 9355 19839
rect 9413 19805 9447 19839
rect 9597 19805 9631 19839
rect 11437 19805 11471 19839
rect 14841 19805 14875 19839
rect 14933 19805 14967 19839
rect 15485 19805 15519 19839
rect 15577 19805 15611 19839
rect 15761 19805 15795 19839
rect 16129 19805 16163 19839
rect 16497 19805 16531 19839
rect 18245 19805 18279 19839
rect 19993 19805 20027 19839
rect 21833 19805 21867 19839
rect 24593 19805 24627 19839
rect 25237 19805 25271 19839
rect 2053 19737 2087 19771
rect 8401 19737 8435 19771
rect 11805 19737 11839 19771
rect 16589 19737 16623 19771
rect 16789 19737 16823 19771
rect 20545 19737 20579 19771
rect 21097 19737 21131 19771
rect 23857 19737 23891 19771
rect 23949 19737 23983 19771
rect 3525 19669 3559 19703
rect 4261 19669 4295 19703
rect 5089 19669 5123 19703
rect 6469 19669 6503 19703
rect 11253 19669 11287 19703
rect 15301 19669 15335 19703
rect 16129 19669 16163 19703
rect 16957 19669 16991 19703
rect 18061 19669 18095 19703
rect 18981 19669 19015 19703
rect 19809 19669 19843 19703
rect 21005 19669 21039 19703
rect 21649 19669 21683 19703
rect 23489 19669 23523 19703
rect 24409 19669 24443 19703
rect 1593 19465 1627 19499
rect 2421 19465 2455 19499
rect 6929 19465 6963 19499
rect 9413 19465 9447 19499
rect 10977 19465 11011 19499
rect 12357 19465 12391 19499
rect 13277 19465 13311 19499
rect 21373 19465 21407 19499
rect 25237 19465 25271 19499
rect 6561 19397 6595 19431
rect 7941 19397 7975 19431
rect 12817 19397 12851 19431
rect 14565 19397 14599 19431
rect 18061 19397 18095 19431
rect 22201 19397 22235 19431
rect 23765 19397 23799 19431
rect 1501 19329 1535 19363
rect 1961 19329 1995 19363
rect 2605 19329 2639 19363
rect 2697 19329 2731 19363
rect 5089 19329 5123 19363
rect 5273 19329 5307 19363
rect 5365 19329 5399 19363
rect 5549 19329 5583 19363
rect 6469 19329 6503 19363
rect 6653 19329 6687 19363
rect 6837 19329 6871 19363
rect 7021 19329 7055 19363
rect 7665 19329 7699 19363
rect 13093 19329 13127 19363
rect 15301 19329 15335 19363
rect 16037 19329 16071 19363
rect 16221 19329 16255 19363
rect 16313 19329 16347 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17785 19329 17819 19363
rect 21649 19329 21683 19363
rect 23397 19329 23431 19363
rect 23489 19329 23523 19363
rect 2973 19261 3007 19295
rect 4445 19261 4479 19295
rect 11069 19261 11103 19295
rect 11253 19261 11287 19295
rect 12449 19261 12483 19295
rect 12633 19261 12667 19295
rect 12909 19261 12943 19295
rect 14933 19261 14967 19295
rect 15025 19261 15059 19295
rect 15761 19261 15795 19295
rect 19625 19261 19659 19295
rect 19901 19261 19935 19295
rect 15853 19193 15887 19227
rect 21465 19193 21499 19227
rect 22385 19193 22419 19227
rect 2145 19125 2179 19159
rect 4905 19125 4939 19159
rect 5825 19125 5859 19159
rect 10609 19125 10643 19159
rect 11989 19125 12023 19159
rect 13093 19125 13127 19159
rect 15209 19125 15243 19159
rect 15485 19125 15519 19159
rect 16773 19125 16807 19159
rect 19533 19125 19567 19159
rect 23213 19125 23247 19159
rect 3801 18921 3835 18955
rect 6469 18921 6503 18955
rect 8493 18921 8527 18955
rect 11621 18921 11655 18955
rect 14197 18921 14231 18955
rect 14565 18921 14599 18955
rect 15393 18921 15427 18955
rect 15853 18921 15887 18955
rect 16037 18921 16071 18955
rect 16497 18921 16531 18955
rect 18153 18921 18187 18955
rect 19533 18921 19567 18955
rect 24869 18921 24903 18955
rect 25421 18921 25455 18955
rect 5641 18853 5675 18887
rect 8309 18853 8343 18887
rect 15577 18853 15611 18887
rect 17785 18853 17819 18887
rect 19257 18853 19291 18887
rect 24685 18853 24719 18887
rect 4353 18785 4387 18819
rect 9873 18785 9907 18819
rect 14933 18785 14967 18819
rect 15850 18785 15884 18819
rect 16221 18785 16255 18819
rect 17877 18785 17911 18819
rect 18797 18785 18831 18819
rect 20637 18785 20671 18819
rect 24409 18785 24443 18819
rect 4261 18717 4295 18751
rect 4721 18717 4755 18751
rect 4905 18717 4939 18751
rect 5089 18717 5123 18751
rect 5917 18717 5951 18751
rect 11989 18717 12023 18751
rect 14105 18717 14139 18751
rect 14657 18717 14691 18751
rect 14841 18717 14875 18751
rect 15025 18717 15059 18751
rect 15209 18717 15243 18751
rect 15485 18717 15519 18751
rect 15761 18717 15795 18751
rect 16313 18717 16347 18751
rect 16589 18717 16623 18751
rect 16957 18717 16991 18751
rect 17141 18717 17175 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 19441 18717 19475 18751
rect 19717 18717 19751 18751
rect 25145 18717 25179 18751
rect 25237 18717 25271 18751
rect 4169 18649 4203 18683
rect 8033 18649 8067 18683
rect 10149 18649 10183 18683
rect 16037 18649 16071 18683
rect 17417 18649 17451 18683
rect 20913 18649 20947 18683
rect 4813 18581 4847 18615
rect 11805 18581 11839 18615
rect 16681 18581 16715 18615
rect 17325 18581 17359 18615
rect 22385 18581 22419 18615
rect 24961 18581 24995 18615
rect 8953 18377 8987 18411
rect 10333 18377 10367 18411
rect 13277 18377 13311 18411
rect 14105 18377 14139 18411
rect 21833 18377 21867 18411
rect 22293 18377 22327 18411
rect 4629 18309 4663 18343
rect 7297 18309 7331 18343
rect 15393 18309 15427 18343
rect 16313 18309 16347 18343
rect 18245 18309 18279 18343
rect 22201 18309 22235 18343
rect 23397 18309 23431 18343
rect 1501 18241 1535 18275
rect 2329 18241 2363 18275
rect 7021 18241 7055 18275
rect 7481 18241 7515 18275
rect 7665 18241 7699 18275
rect 7757 18241 7791 18275
rect 8585 18241 8619 18275
rect 10149 18241 10183 18275
rect 10517 18241 10551 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 14381 18241 14415 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 16037 18241 16071 18275
rect 16681 18241 16715 18275
rect 17141 18241 17175 18275
rect 17693 18241 17727 18275
rect 17877 18241 17911 18275
rect 19993 18241 20027 18275
rect 21465 18241 21499 18275
rect 25513 18241 25547 18275
rect 4353 18173 4387 18207
rect 7297 18173 7331 18207
rect 8033 18173 8067 18207
rect 8493 18173 8527 18207
rect 9505 18173 9539 18207
rect 11529 18173 11563 18207
rect 11805 18173 11839 18207
rect 16773 18173 16807 18207
rect 17417 18173 17451 18207
rect 18061 18173 18095 18207
rect 22385 18173 22419 18207
rect 23121 18173 23155 18207
rect 7481 18105 7515 18139
rect 15945 18105 15979 18139
rect 1593 18037 1627 18071
rect 2145 18037 2179 18071
rect 6101 18037 6135 18071
rect 7113 18037 7147 18071
rect 8125 18037 8159 18071
rect 8309 18037 8343 18071
rect 16681 18037 16715 18071
rect 17049 18037 17083 18071
rect 17233 18037 17267 18071
rect 17325 18037 17359 18071
rect 21281 18037 21315 18071
rect 24869 18037 24903 18071
rect 25329 18037 25363 18071
rect 6745 17833 6779 17867
rect 9045 17833 9079 17867
rect 9965 17833 9999 17867
rect 10609 17833 10643 17867
rect 11989 17833 12023 17867
rect 15669 17833 15703 17867
rect 19257 17833 19291 17867
rect 23121 17833 23155 17867
rect 24133 17833 24167 17867
rect 8677 17765 8711 17799
rect 9781 17765 9815 17799
rect 23581 17765 23615 17799
rect 23949 17765 23983 17799
rect 24409 17765 24443 17799
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 3433 17697 3467 17731
rect 4261 17697 4295 17731
rect 9413 17697 9447 17731
rect 11805 17697 11839 17731
rect 14657 17697 14691 17731
rect 16037 17697 16071 17731
rect 19901 17697 19935 17731
rect 23213 17697 23247 17731
rect 23673 17697 23707 17731
rect 24869 17697 24903 17731
rect 24961 17697 24995 17731
rect 3985 17629 4019 17663
rect 4169 17629 4203 17663
rect 5273 17629 5307 17663
rect 7389 17629 7423 17663
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 8125 17629 8159 17663
rect 8493 17629 8527 17663
rect 8585 17629 8619 17663
rect 8769 17629 8803 17663
rect 8953 17629 8987 17663
rect 10793 17629 10827 17663
rect 11989 17629 12023 17663
rect 15577 17629 15611 17663
rect 15853 17629 15887 17663
rect 15945 17629 15979 17663
rect 16221 17629 16255 17663
rect 20545 17629 20579 17663
rect 22385 17629 22419 17663
rect 23121 17629 23155 17663
rect 23397 17629 23431 17663
rect 24777 17629 24811 17663
rect 9505 17561 9539 17595
rect 11713 17561 11747 17595
rect 15485 17561 15519 17595
rect 19717 17561 19751 17595
rect 20821 17561 20855 17595
rect 3801 17493 3835 17527
rect 8493 17493 8527 17527
rect 12173 17493 12207 17527
rect 16129 17493 16163 17527
rect 19625 17493 19659 17527
rect 22293 17493 22327 17527
rect 23029 17493 23063 17527
rect 2237 17289 2271 17323
rect 3065 17289 3099 17323
rect 4077 17289 4111 17323
rect 6653 17289 6687 17323
rect 7389 17289 7423 17323
rect 9137 17289 9171 17323
rect 10885 17289 10919 17323
rect 16957 17289 16991 17323
rect 21097 17289 21131 17323
rect 22293 17289 22327 17323
rect 25329 17289 25363 17323
rect 4629 17221 4663 17255
rect 8401 17221 8435 17255
rect 11897 17221 11931 17255
rect 11989 17221 12023 17255
rect 22201 17221 22235 17255
rect 23857 17221 23891 17255
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 2421 17153 2455 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 3709 17153 3743 17187
rect 3893 17153 3927 17187
rect 4353 17153 4387 17187
rect 6377 17153 6411 17187
rect 6929 17153 6963 17187
rect 7665 17153 7699 17187
rect 8135 17153 8169 17187
rect 8677 17153 8711 17187
rect 11069 17153 11103 17187
rect 11345 17153 11379 17187
rect 12541 17153 12575 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 16681 17153 16715 17187
rect 19625 17153 19659 17187
rect 19809 17153 19843 17187
rect 20637 17153 20671 17187
rect 21281 17153 21315 17187
rect 23581 17153 23615 17187
rect 25053 17153 25087 17187
rect 25513 17153 25547 17187
rect 3157 17085 3191 17119
rect 6101 17085 6135 17119
rect 6653 17085 6687 17119
rect 7757 17085 7791 17119
rect 12081 17085 12115 17119
rect 12817 17085 12851 17119
rect 16957 17085 16991 17119
rect 20729 17085 20763 17119
rect 22385 17085 22419 17119
rect 1593 17017 1627 17051
rect 3525 17017 3559 17051
rect 3617 17017 3651 17051
rect 8033 17017 8067 17051
rect 11529 17017 11563 17051
rect 13369 17017 13403 17051
rect 15945 17017 15979 17051
rect 21833 17017 21867 17051
rect 24133 17017 24167 17051
rect 25237 17017 25271 17051
rect 1869 16949 1903 16983
rect 2605 16949 2639 16983
rect 3893 16949 3927 16983
rect 6469 16949 6503 16983
rect 7205 16949 7239 16983
rect 8769 16949 8803 16983
rect 11161 16949 11195 16983
rect 12357 16949 12391 16983
rect 14933 16949 14967 16983
rect 15301 16949 15335 16983
rect 15669 16949 15703 16983
rect 16773 16949 16807 16983
rect 19625 16949 19659 16983
rect 20913 16949 20947 16983
rect 23397 16949 23431 16983
rect 24317 16949 24351 16983
rect 6009 16745 6043 16779
rect 6377 16745 6411 16779
rect 10425 16745 10459 16779
rect 11326 16745 11360 16779
rect 19901 16745 19935 16779
rect 21741 16745 21775 16779
rect 22109 16745 22143 16779
rect 4537 16677 4571 16711
rect 5273 16677 5307 16711
rect 5825 16677 5859 16711
rect 10333 16677 10367 16711
rect 10793 16677 10827 16711
rect 18797 16677 18831 16711
rect 19993 16677 20027 16711
rect 22477 16677 22511 16711
rect 1593 16609 1627 16643
rect 1869 16609 1903 16643
rect 3341 16609 3375 16643
rect 3801 16609 3835 16643
rect 4905 16609 4939 16643
rect 13737 16609 13771 16643
rect 14749 16609 14783 16643
rect 15393 16609 15427 16643
rect 15669 16609 15703 16643
rect 17877 16609 17911 16643
rect 18245 16609 18279 16643
rect 19257 16609 19291 16643
rect 20453 16609 20487 16643
rect 20637 16609 20671 16643
rect 20821 16609 20855 16643
rect 21373 16609 21407 16643
rect 24501 16609 24535 16643
rect 3617 16541 3651 16575
rect 4813 16541 4847 16575
rect 6193 16541 6227 16575
rect 6561 16541 6595 16575
rect 8125 16541 8159 16575
rect 8217 16541 8251 16575
rect 8309 16541 8343 16575
rect 8493 16541 8527 16575
rect 8585 16541 8619 16575
rect 8769 16541 8803 16575
rect 11069 16541 11103 16575
rect 14657 16541 14691 16575
rect 15301 16541 15335 16575
rect 16221 16541 16255 16575
rect 18061 16541 18095 16575
rect 18337 16541 18371 16575
rect 18429 16541 18463 16575
rect 19073 16541 19107 16575
rect 21005 16541 21039 16575
rect 21465 16541 21499 16575
rect 22006 16543 22040 16577
rect 23765 16541 23799 16575
rect 24041 16541 24075 16575
rect 25329 16541 25363 16575
rect 4537 16473 4571 16507
rect 5457 16473 5491 16507
rect 8677 16473 8711 16507
rect 9965 16473 9999 16507
rect 10517 16473 10551 16507
rect 13553 16473 13587 16507
rect 16773 16473 16807 16507
rect 18797 16473 18831 16507
rect 3433 16405 3467 16439
rect 4445 16405 4479 16439
rect 4721 16405 4755 16439
rect 5365 16405 5399 16439
rect 5917 16405 5951 16439
rect 7849 16405 7883 16439
rect 10977 16405 11011 16439
rect 12817 16405 12851 16439
rect 13185 16405 13219 16439
rect 13645 16405 13679 16439
rect 15025 16405 15059 16439
rect 18981 16405 19015 16439
rect 20361 16405 20395 16439
rect 21005 16405 21039 16439
rect 21925 16405 21959 16439
rect 23581 16405 23615 16439
rect 23857 16405 23891 16439
rect 25053 16405 25087 16439
rect 25145 16405 25179 16439
rect 3065 16201 3099 16235
rect 4261 16201 4295 16235
rect 9689 16201 9723 16235
rect 10425 16201 10459 16235
rect 12265 16201 12299 16235
rect 15761 16201 15795 16235
rect 18981 16201 19015 16235
rect 19625 16201 19659 16235
rect 22293 16201 22327 16235
rect 22845 16201 22879 16235
rect 23305 16201 23339 16235
rect 25421 16201 25455 16235
rect 3157 16133 3191 16167
rect 3341 16133 3375 16167
rect 8217 16133 8251 16167
rect 15669 16133 15703 16167
rect 21097 16133 21131 16167
rect 21833 16133 21867 16167
rect 23949 16133 23983 16167
rect 1501 16065 1535 16099
rect 4169 16065 4203 16099
rect 4353 16065 4387 16099
rect 5917 16065 5951 16099
rect 7941 16065 7975 16099
rect 10517 16065 10551 16099
rect 11805 16065 11839 16099
rect 11989 16065 12023 16099
rect 12081 16065 12115 16099
rect 17141 16065 17175 16099
rect 19165 16065 19199 16099
rect 19717 16065 19751 16099
rect 21005 16065 21039 16099
rect 23213 16065 23247 16099
rect 2605 15997 2639 16031
rect 3525 15997 3559 16031
rect 9965 15997 9999 16031
rect 10885 15997 10919 16031
rect 12449 15997 12483 16031
rect 12725 15997 12759 16031
rect 15853 15997 15887 16031
rect 17233 15997 17267 16031
rect 17509 15997 17543 16031
rect 21189 15997 21223 16031
rect 23397 15997 23431 16031
rect 23673 15997 23707 16031
rect 2881 15929 2915 15963
rect 10333 15929 10367 15963
rect 11161 15929 11195 15963
rect 16957 15929 16991 15963
rect 22201 15929 22235 15963
rect 1593 15861 1627 15895
rect 2237 15861 2271 15895
rect 5733 15861 5767 15895
rect 10701 15861 10735 15895
rect 11345 15861 11379 15895
rect 12081 15861 12115 15895
rect 14197 15861 14231 15895
rect 15301 15861 15335 15895
rect 19441 15861 19475 15895
rect 20361 15861 20395 15895
rect 20637 15861 20671 15895
rect 9413 15657 9447 15691
rect 11621 15657 11655 15691
rect 12541 15657 12575 15691
rect 12909 15657 12943 15691
rect 19520 15657 19554 15691
rect 21005 15657 21039 15691
rect 24409 15657 24443 15691
rect 25421 15657 25455 15691
rect 18889 15589 18923 15623
rect 4997 15521 5031 15555
rect 14933 15521 14967 15555
rect 15945 15521 15979 15555
rect 19257 15521 19291 15555
rect 22477 15521 22511 15555
rect 24869 15521 24903 15555
rect 24961 15521 24995 15555
rect 2697 15453 2731 15487
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 3065 15453 3099 15487
rect 3249 15453 3283 15487
rect 3801 15453 3835 15487
rect 4629 15453 4663 15487
rect 4813 15453 4847 15487
rect 7021 15453 7055 15487
rect 8217 15453 8251 15487
rect 8493 15453 8527 15487
rect 9597 15453 9631 15487
rect 10333 15453 10367 15487
rect 11069 15453 11103 15487
rect 11437 15453 11471 15487
rect 12725 15453 12759 15487
rect 13093 15453 13127 15487
rect 15117 15453 15151 15487
rect 18061 15453 18095 15487
rect 18705 15453 18739 15487
rect 22385 15453 22419 15487
rect 25237 15453 25271 15487
rect 4445 15385 4479 15419
rect 4721 15385 4755 15419
rect 5273 15385 5307 15419
rect 16221 15385 16255 15419
rect 17969 15385 18003 15419
rect 18337 15385 18371 15419
rect 22753 15385 22787 15419
rect 24777 15385 24811 15419
rect 2513 15317 2547 15351
rect 3157 15317 3191 15351
rect 10517 15317 10551 15351
rect 11253 15317 11287 15351
rect 15301 15317 15335 15351
rect 22201 15317 22235 15351
rect 24225 15317 24259 15351
rect 5733 15113 5767 15147
rect 9965 15113 9999 15147
rect 18245 15113 18279 15147
rect 19165 15113 19199 15147
rect 19809 15113 19843 15147
rect 22385 15113 22419 15147
rect 22937 15113 22971 15147
rect 24869 15113 24903 15147
rect 3433 15045 3467 15079
rect 3617 15045 3651 15079
rect 13093 15045 13127 15079
rect 18889 15045 18923 15079
rect 1593 14977 1627 15011
rect 4169 14977 4203 15011
rect 5273 14977 5307 15011
rect 6561 14977 6595 15011
rect 7205 14977 7239 15011
rect 11713 14977 11747 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 15369 14977 15403 15011
rect 18429 14977 18463 15011
rect 18613 14977 18647 15011
rect 19441 14977 19475 15011
rect 19993 14977 20027 15011
rect 20821 14977 20855 15011
rect 22293 14977 22327 15011
rect 23121 14977 23155 15011
rect 24961 14977 24995 15011
rect 1869 14909 1903 14943
rect 3801 14909 3835 14943
rect 7297 14909 7331 14943
rect 7481 14909 7515 14943
rect 9505 14909 9539 14943
rect 10793 14909 10827 14943
rect 11253 14909 11287 14943
rect 15025 14909 15059 14943
rect 17693 14909 17727 14943
rect 18153 14909 18187 14943
rect 19349 14909 19383 14943
rect 19533 14909 19567 14943
rect 19625 14909 19659 14943
rect 22477 14909 22511 14943
rect 23397 14909 23431 14943
rect 3341 14841 3375 14875
rect 4537 14841 4571 14875
rect 5549 14841 5583 14875
rect 6837 14841 6871 14875
rect 9873 14841 9907 14875
rect 11069 14841 11103 14875
rect 14381 14841 14415 14875
rect 15209 14841 15243 14875
rect 18061 14841 18095 14875
rect 25237 14841 25271 14875
rect 4629 14773 4663 14807
rect 6377 14773 6411 14807
rect 11529 14773 11563 14807
rect 20637 14773 20671 14807
rect 21925 14773 21959 14807
rect 25421 14773 25455 14807
rect 2237 14569 2271 14603
rect 3065 14569 3099 14603
rect 13829 14569 13863 14603
rect 18705 14569 18739 14603
rect 22477 14569 22511 14603
rect 24041 14569 24075 14603
rect 24961 14569 24995 14603
rect 25421 14569 25455 14603
rect 2881 14501 2915 14535
rect 5365 14501 5399 14535
rect 9689 14501 9723 14535
rect 18521 14501 18555 14535
rect 23949 14501 23983 14535
rect 24685 14501 24719 14535
rect 2973 14433 3007 14467
rect 5825 14433 5859 14467
rect 14841 14433 14875 14467
rect 16589 14433 16623 14467
rect 20729 14433 20763 14467
rect 1409 14365 1443 14399
rect 2421 14365 2455 14399
rect 2513 14365 2547 14399
rect 3249 14365 3283 14399
rect 5549 14365 5583 14399
rect 8033 14365 8067 14399
rect 9873 14365 9907 14399
rect 10609 14365 10643 14399
rect 14565 14365 14599 14399
rect 16773 14365 16807 14399
rect 20453 14365 20487 14399
rect 22661 14365 22695 14399
rect 24501 14365 24535 14399
rect 25145 14365 25179 14399
rect 25237 14365 25271 14399
rect 4997 14297 5031 14331
rect 8309 14297 8343 14331
rect 10885 14297 10919 14331
rect 13553 14297 13587 14331
rect 18245 14297 18279 14331
rect 23581 14297 23615 14331
rect 1593 14229 1627 14263
rect 5457 14229 5491 14263
rect 7297 14229 7331 14263
rect 12357 14229 12391 14263
rect 16865 14229 16899 14263
rect 22201 14229 22235 14263
rect 1593 14025 1627 14059
rect 3157 14025 3191 14059
rect 3525 14025 3559 14059
rect 6377 14025 6411 14059
rect 10793 14025 10827 14059
rect 10885 14025 10919 14059
rect 11529 14025 11563 14059
rect 11897 14025 11931 14059
rect 11989 14025 12023 14059
rect 15577 14025 15611 14059
rect 15945 14025 15979 14059
rect 21465 14025 21499 14059
rect 24041 13957 24075 13991
rect 1409 13889 1443 13923
rect 3065 13889 3099 13923
rect 3617 13889 3651 13923
rect 5641 13889 5675 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 8493 13889 8527 13923
rect 11069 13889 11103 13923
rect 12541 13889 12575 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 14749 13889 14783 13923
rect 14933 13889 14967 13923
rect 15761 13889 15795 13923
rect 16129 13889 16163 13923
rect 17693 13889 17727 13923
rect 3801 13821 3835 13855
rect 4905 13821 4939 13855
rect 6929 13821 6963 13855
rect 8769 13821 8803 13855
rect 10241 13821 10275 13855
rect 10333 13821 10367 13855
rect 12081 13821 12115 13855
rect 15025 13821 15059 13855
rect 15485 13821 15519 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 23765 13821 23799 13855
rect 25513 13821 25547 13855
rect 5273 13753 5307 13787
rect 10701 13753 10735 13787
rect 15301 13753 15335 13787
rect 2881 13685 2915 13719
rect 5365 13685 5399 13719
rect 5457 13685 5491 13719
rect 8401 13685 8435 13719
rect 12357 13685 12391 13719
rect 14289 13685 14323 13719
rect 17509 13685 17543 13719
rect 6653 13481 6687 13515
rect 9045 13481 9079 13515
rect 11161 13481 11195 13515
rect 13829 13481 13863 13515
rect 18153 13481 18187 13515
rect 19901 13481 19935 13515
rect 21005 13481 21039 13515
rect 21373 13481 21407 13515
rect 24501 13481 24535 13515
rect 25145 13481 25179 13515
rect 7205 13413 7239 13447
rect 20177 13413 20211 13447
rect 4353 13345 4387 13379
rect 6929 13345 6963 13379
rect 7389 13345 7423 13379
rect 8125 13345 8159 13379
rect 9873 13345 9907 13379
rect 9965 13345 9999 13379
rect 11805 13345 11839 13379
rect 16405 13345 16439 13379
rect 20729 13345 20763 13379
rect 3341 13277 3375 13311
rect 4813 13277 4847 13311
rect 6837 13277 6871 13311
rect 8033 13277 8067 13311
rect 9229 13277 9263 13311
rect 12081 13277 12115 13311
rect 14105 13277 14139 13311
rect 16313 13277 16347 13311
rect 18245 13277 18279 13311
rect 18613 13277 18647 13311
rect 19441 13277 19475 13311
rect 20085 13277 20119 13311
rect 21189 13277 21223 13311
rect 21557 13277 21591 13311
rect 23949 13277 23983 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25237 13277 25271 13311
rect 1501 13209 1535 13243
rect 4169 13209 4203 13243
rect 7941 13209 7975 13243
rect 11529 13209 11563 13243
rect 12357 13209 12391 13243
rect 14381 13209 14415 13243
rect 16681 13209 16715 13243
rect 20545 13209 20579 13243
rect 1593 13141 1627 13175
rect 3157 13141 3191 13175
rect 3801 13141 3835 13175
rect 4261 13141 4295 13175
rect 4629 13141 4663 13175
rect 7573 13141 7607 13175
rect 9413 13141 9447 13175
rect 9781 13141 9815 13175
rect 11621 13141 11655 13175
rect 15853 13141 15887 13175
rect 16129 13141 16163 13175
rect 18429 13141 18463 13175
rect 18797 13141 18831 13175
rect 19257 13141 19291 13175
rect 20637 13141 20671 13175
rect 23765 13141 23799 13175
rect 25421 13141 25455 13175
rect 4537 12937 4571 12971
rect 7205 12937 7239 12971
rect 8493 12937 8527 12971
rect 13277 12937 13311 12971
rect 13461 12937 13495 12971
rect 15025 12937 15059 12971
rect 16681 12937 16715 12971
rect 17969 12937 18003 12971
rect 20913 12937 20947 12971
rect 21465 12937 21499 12971
rect 24409 12937 24443 12971
rect 25053 12937 25087 12971
rect 3065 12869 3099 12903
rect 14013 12869 14047 12903
rect 14565 12869 14599 12903
rect 15209 12869 15243 12903
rect 15577 12869 15611 12903
rect 17049 12869 17083 12903
rect 17509 12869 17543 12903
rect 24593 12869 24627 12903
rect 2421 12801 2455 12835
rect 4905 12801 4939 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 7849 12801 7883 12835
rect 8217 12801 8251 12835
rect 10425 12801 10459 12835
rect 10701 12801 10735 12835
rect 11069 12801 11103 12835
rect 11897 12801 11931 12835
rect 12449 12801 12483 12835
rect 13093 12801 13127 12835
rect 13645 12801 13679 12835
rect 18061 12801 18095 12835
rect 20085 12801 20119 12835
rect 22661 12801 22695 12835
rect 25329 12801 25363 12835
rect 2789 12733 2823 12767
rect 7665 12733 7699 12767
rect 10517 12733 10551 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 14473 12733 14507 12767
rect 17141 12733 17175 12767
rect 17325 12733 17359 12767
rect 18337 12733 18371 12767
rect 19809 12733 19843 12767
rect 20453 12733 20487 12767
rect 21005 12733 21039 12767
rect 22937 12733 22971 12767
rect 13001 12665 13035 12699
rect 14289 12665 14323 12699
rect 14841 12665 14875 12699
rect 17785 12665 17819 12699
rect 20269 12665 20303 12699
rect 20729 12665 20763 12699
rect 21281 12665 21315 12699
rect 24869 12665 24903 12699
rect 25513 12665 25547 12699
rect 2237 12597 2271 12631
rect 4721 12597 4755 12631
rect 7849 12597 7883 12631
rect 8033 12597 8067 12631
rect 10701 12597 10735 12631
rect 10885 12597 10919 12631
rect 11253 12597 11287 12631
rect 11529 12597 11563 12631
rect 3157 12393 3191 12427
rect 5733 12393 5767 12427
rect 12633 12393 12667 12427
rect 13461 12393 13495 12427
rect 14749 12393 14783 12427
rect 18245 12393 18279 12427
rect 19073 12393 19107 12427
rect 19533 12393 19567 12427
rect 23857 12393 23891 12427
rect 12725 12325 12759 12359
rect 13277 12325 13311 12359
rect 17049 12325 17083 12359
rect 18889 12325 18923 12359
rect 22293 12325 22327 12359
rect 23765 12325 23799 12359
rect 3893 12257 3927 12291
rect 4169 12257 4203 12291
rect 6377 12257 6411 12291
rect 10149 12257 10183 12291
rect 11161 12257 11195 12291
rect 17601 12257 17635 12291
rect 18613 12257 18647 12291
rect 20545 12257 20579 12291
rect 1409 12189 1443 12223
rect 6101 12189 6135 12223
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 7757 12189 7791 12223
rect 9965 12189 9999 12223
rect 10885 12189 10919 12223
rect 12909 12189 12943 12223
rect 13553 12189 13587 12223
rect 13645 12189 13679 12223
rect 13737 12189 13771 12223
rect 14933 12189 14967 12223
rect 17509 12189 17543 12223
rect 17877 12189 17911 12223
rect 18429 12189 18463 12223
rect 19441 12189 19475 12223
rect 20453 12189 20487 12223
rect 23397 12189 23431 12223
rect 1685 12121 1719 12155
rect 13001 12121 13035 12155
rect 20821 12121 20855 12155
rect 5641 12053 5675 12087
rect 6193 12053 6227 12087
rect 7113 12053 7147 12087
rect 9597 12053 9631 12087
rect 10057 12053 10091 12087
rect 17417 12053 17451 12087
rect 18061 12053 18095 12087
rect 20269 12053 20303 12087
rect 2421 11849 2455 11883
rect 4537 11849 4571 11883
rect 4629 11849 4663 11883
rect 7481 11849 7515 11883
rect 8401 11849 8435 11883
rect 11345 11849 11379 11883
rect 21465 11849 21499 11883
rect 21833 11849 21867 11883
rect 24869 11849 24903 11883
rect 3065 11781 3099 11815
rect 10885 11781 10919 11815
rect 22201 11781 22235 11815
rect 1409 11713 1443 11747
rect 4813 11713 4847 11747
rect 6561 11713 6595 11747
rect 6745 11713 6779 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 8125 11713 8159 11747
rect 9597 11713 9631 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 12265 11713 12299 11747
rect 15393 11713 15427 11747
rect 15577 11713 15611 11747
rect 17325 11713 17359 11747
rect 20913 11713 20947 11747
rect 21649 11713 21683 11747
rect 24777 11713 24811 11747
rect 1961 11645 1995 11679
rect 2789 11645 2823 11679
rect 4905 11645 4939 11679
rect 5365 11645 5399 11679
rect 11069 11645 11103 11679
rect 11989 11645 12023 11679
rect 21373 11645 21407 11679
rect 22293 11645 22327 11679
rect 22385 11645 22419 11679
rect 24961 11645 24995 11679
rect 2329 11577 2363 11611
rect 5181 11577 5215 11611
rect 11805 11577 11839 11611
rect 12081 11577 12115 11611
rect 21189 11577 21223 11611
rect 1593 11509 1627 11543
rect 6653 11509 6687 11543
rect 9413 11509 9447 11543
rect 10885 11509 10919 11543
rect 15485 11509 15519 11543
rect 17509 11509 17543 11543
rect 24409 11509 24443 11543
rect 4445 11305 4479 11339
rect 4997 11305 5031 11339
rect 6745 11305 6779 11339
rect 7205 11305 7239 11339
rect 9400 11305 9434 11339
rect 10885 11305 10919 11339
rect 14565 11305 14599 11339
rect 15485 11305 15519 11339
rect 17785 11305 17819 11339
rect 22845 11305 22879 11339
rect 25329 11305 25363 11339
rect 7389 11237 7423 11271
rect 8309 11237 8343 11271
rect 15301 11237 15335 11271
rect 17693 11237 17727 11271
rect 18153 11237 18187 11271
rect 20269 11237 20303 11271
rect 24041 11237 24075 11271
rect 3065 11169 3099 11203
rect 6561 11169 6595 11203
rect 15025 11169 15059 11203
rect 16037 11169 16071 11203
rect 16129 11169 16163 11203
rect 17877 11169 17911 11203
rect 18337 11169 18371 11203
rect 20821 11169 20855 11203
rect 23673 11169 23707 11203
rect 24133 11169 24167 11203
rect 4353 11101 4387 11135
rect 4905 11101 4939 11135
rect 5457 11101 5491 11135
rect 5641 11101 5675 11135
rect 6469 11101 6503 11135
rect 6929 11101 6963 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 11253 11101 11287 11135
rect 14473 11101 14507 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 16313 11101 16347 11135
rect 18613 11101 18647 11135
rect 20637 11101 20671 11135
rect 21281 11101 21315 11135
rect 23029 11101 23063 11135
rect 24593 11101 24627 11135
rect 24869 11101 24903 11135
rect 25513 11101 25547 11135
rect 1501 11033 1535 11067
rect 3617 11033 3651 11067
rect 17325 11033 17359 11067
rect 20729 11033 20763 11067
rect 1593 10965 1627 10999
rect 4813 10965 4847 10999
rect 5365 10965 5399 10999
rect 5549 10965 5583 10999
rect 8401 10965 8435 10999
rect 11069 10965 11103 10999
rect 14933 10965 14967 10999
rect 16497 10965 16531 10999
rect 18429 10965 18463 10999
rect 21097 10965 21131 10999
rect 24409 10965 24443 10999
rect 24685 10965 24719 10999
rect 9413 10761 9447 10795
rect 10885 10761 10919 10795
rect 12633 10761 12667 10795
rect 18613 10761 18647 10795
rect 18797 10761 18831 10795
rect 21833 10761 21867 10795
rect 6009 10693 6043 10727
rect 12725 10693 12759 10727
rect 12909 10693 12943 10727
rect 20085 10693 20119 10727
rect 23581 10693 23615 10727
rect 1501 10625 1535 10659
rect 2697 10625 2731 10659
rect 4537 10625 4571 10659
rect 4629 10625 4663 10659
rect 4721 10625 4755 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 5365 10625 5399 10659
rect 5733 10625 5767 10659
rect 6745 10625 6779 10659
rect 9597 10625 9631 10659
rect 13645 10625 13679 10659
rect 14473 10625 14507 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16037 10625 16071 10659
rect 16221 10625 16255 10659
rect 16865 10625 16899 10659
rect 18981 10625 19015 10659
rect 22017 10625 22051 10659
rect 23305 10625 23339 10659
rect 25237 10625 25271 10659
rect 1961 10557 1995 10591
rect 2421 10557 2455 10591
rect 5457 10557 5491 10591
rect 6009 10557 6043 10591
rect 7665 10557 7699 10591
rect 7941 10557 7975 10591
rect 12173 10557 12207 10591
rect 14749 10557 14783 10591
rect 15301 10557 15335 10591
rect 15577 10557 15611 10591
rect 17141 10557 17175 10591
rect 19809 10557 19843 10591
rect 22753 10557 22787 10591
rect 2329 10489 2363 10523
rect 5825 10489 5859 10523
rect 7205 10489 7239 10523
rect 12541 10489 12575 10523
rect 23121 10489 23155 10523
rect 1593 10421 1627 10455
rect 2513 10421 2547 10455
rect 4261 10421 4295 10455
rect 5641 10421 5675 10455
rect 6929 10421 6963 10455
rect 13093 10421 13127 10455
rect 13737 10421 13771 10455
rect 14105 10421 14139 10455
rect 21557 10421 21591 10455
rect 23213 10421 23247 10455
rect 25053 10421 25087 10455
rect 25421 10421 25455 10455
rect 5457 10217 5491 10251
rect 7389 10217 7423 10251
rect 8401 10217 8435 10251
rect 10333 10217 10367 10251
rect 12081 10217 12115 10251
rect 15945 10217 15979 10251
rect 16681 10217 16715 10251
rect 20821 10217 20855 10251
rect 22845 10217 22879 10251
rect 10241 10149 10275 10183
rect 11989 10149 12023 10183
rect 14197 10149 14231 10183
rect 15025 10149 15059 10183
rect 20637 10149 20671 10183
rect 24685 10149 24719 10183
rect 1409 10081 1443 10115
rect 1685 10081 1719 10115
rect 5181 10081 5215 10115
rect 9873 10081 9907 10115
rect 11621 10081 11655 10115
rect 12449 10081 12483 10115
rect 12817 10081 12851 10115
rect 13369 10081 13403 10115
rect 14749 10081 14783 10115
rect 15209 10081 15243 10115
rect 17325 10081 17359 10115
rect 19901 10081 19935 10115
rect 20361 10081 20395 10115
rect 21465 10081 21499 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 24409 10081 24443 10115
rect 3249 10013 3283 10047
rect 5089 10013 5123 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 8585 10013 8619 10047
rect 9505 10013 9539 10047
rect 10609 10013 10643 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 12357 10013 12391 10047
rect 13001 10013 13035 10047
rect 13461 10013 13495 10047
rect 14381 10013 14415 10047
rect 14565 10013 14599 10047
rect 14657 10007 14691 10041
rect 15669 10013 15703 10047
rect 15761 10013 15795 10047
rect 16405 10013 16439 10047
rect 17049 10013 17083 10047
rect 19625 10013 19659 10047
rect 21281 10013 21315 10047
rect 23857 10013 23891 10047
rect 25145 10013 25179 10047
rect 5641 9945 5675 9979
rect 12633 9945 12667 9979
rect 12725 9945 12759 9979
rect 13737 9945 13771 9979
rect 16037 9945 16071 9979
rect 16219 9945 16253 9979
rect 16497 9945 16531 9979
rect 21373 9945 21407 9979
rect 3157 9877 3191 9911
rect 3341 9877 3375 9911
rect 9321 9877 9355 9911
rect 10425 9877 10459 9911
rect 11437 9877 11471 9911
rect 13277 9877 13311 9911
rect 15301 9877 15335 9911
rect 16697 9877 16731 9911
rect 16865 9877 16899 9911
rect 18797 9877 18831 9911
rect 19257 9877 19291 9911
rect 19717 9877 19751 9911
rect 20913 9877 20947 9911
rect 23213 9877 23247 9911
rect 23673 9877 23707 9911
rect 24869 9877 24903 9911
rect 25421 9877 25455 9911
rect 7941 9673 7975 9707
rect 11529 9673 11563 9707
rect 13001 9673 13035 9707
rect 24961 9673 24995 9707
rect 9045 9605 9079 9639
rect 13093 9605 13127 9639
rect 13293 9605 13327 9639
rect 13737 9605 13771 9639
rect 14749 9605 14783 9639
rect 15393 9605 15427 9639
rect 19993 9605 20027 9639
rect 1501 9537 1535 9571
rect 2789 9537 2823 9571
rect 4169 9537 4203 9571
rect 4261 9537 4295 9571
rect 4445 9537 4479 9571
rect 4537 9537 4571 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 7389 9537 7423 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 8769 9537 8803 9571
rect 11161 9537 11195 9571
rect 11253 9537 11287 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 12449 9537 12483 9571
rect 12550 9537 12584 9571
rect 12817 9537 12851 9571
rect 13553 9537 13587 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14105 9537 14139 9571
rect 14657 9537 14691 9571
rect 15025 9537 15059 9571
rect 15209 9537 15243 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 15853 9537 15887 9571
rect 15945 9537 15979 9571
rect 16129 9537 16163 9571
rect 17601 9537 17635 9571
rect 18245 9537 18279 9571
rect 21465 9537 21499 9571
rect 22661 9537 22695 9571
rect 24869 9537 24903 9571
rect 25513 9537 25547 9571
rect 2697 9469 2731 9503
rect 3341 9469 3375 9503
rect 4905 9469 4939 9503
rect 5181 9469 5215 9503
rect 11897 9469 11931 9503
rect 12633 9469 12667 9503
rect 14289 9469 14323 9503
rect 16773 9469 16807 9503
rect 22937 9469 22971 9503
rect 25053 9469 25087 9503
rect 3617 9401 3651 9435
rect 5273 9401 5307 9435
rect 13461 9401 13495 9435
rect 16037 9401 16071 9435
rect 24409 9401 24443 9435
rect 1593 9333 1627 9367
rect 3065 9333 3099 9367
rect 3801 9333 3835 9367
rect 3985 9333 4019 9367
rect 7665 9333 7699 9367
rect 10517 9333 10551 9367
rect 13277 9333 13311 9367
rect 14197 9333 14231 9367
rect 17325 9333 17359 9367
rect 17877 9333 17911 9367
rect 21281 9333 21315 9367
rect 24501 9333 24535 9367
rect 25329 9333 25363 9367
rect 5733 9129 5767 9163
rect 9689 9129 9723 9163
rect 18889 9129 18923 9163
rect 19698 9129 19732 9163
rect 21189 9129 21223 9163
rect 23305 9129 23339 9163
rect 9505 9061 9539 9095
rect 12265 9061 12299 9095
rect 12357 9061 12391 9095
rect 3249 8993 3283 9027
rect 3525 8993 3559 9027
rect 4261 8993 4295 9027
rect 4353 8993 4387 9027
rect 4997 8993 5031 9027
rect 5641 8993 5675 9027
rect 9229 8993 9263 9027
rect 9781 8993 9815 9027
rect 11437 8993 11471 9027
rect 11897 8993 11931 9027
rect 19441 8993 19475 9027
rect 23673 8993 23707 9027
rect 24961 8993 24995 9027
rect 3157 8925 3191 8959
rect 4169 8925 4203 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 9965 8925 9999 8959
rect 11529 8925 11563 8959
rect 12173 8925 12207 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 13185 8925 13219 8959
rect 13369 8925 13403 8959
rect 16221 8925 16255 8959
rect 17693 8925 17727 8959
rect 18245 8925 18279 8959
rect 19073 8925 19107 8959
rect 21465 8925 21499 8959
rect 23489 8925 23523 8959
rect 25513 8925 25547 8959
rect 24225 8857 24259 8891
rect 24869 8857 24903 8891
rect 3801 8789 3835 8823
rect 5457 8789 5491 8823
rect 5917 8789 5951 8823
rect 10149 8789 10183 8823
rect 11989 8789 12023 8823
rect 12725 8789 12759 8823
rect 16773 8789 16807 8823
rect 17509 8789 17543 8823
rect 18061 8789 18095 8823
rect 21281 8789 21315 8823
rect 24409 8789 24443 8823
rect 24777 8789 24811 8823
rect 25329 8789 25363 8823
rect 5365 8585 5399 8619
rect 9321 8585 9355 8619
rect 14197 8585 14231 8619
rect 15669 8585 15703 8619
rect 15761 8585 15795 8619
rect 17141 8585 17175 8619
rect 19993 8585 20027 8619
rect 20821 8585 20855 8619
rect 21465 8585 21499 8619
rect 9689 8517 9723 8551
rect 9781 8517 9815 8551
rect 12725 8517 12759 8551
rect 20361 8517 20395 8551
rect 21005 8517 21039 8551
rect 24041 8517 24075 8551
rect 1501 8449 1535 8483
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 2513 8449 2547 8483
rect 3718 8449 3752 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4445 8449 4479 8483
rect 4905 8449 4939 8483
rect 7389 8449 7423 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 12173 8449 12207 8483
rect 15209 8449 15243 8483
rect 16957 8449 16991 8483
rect 19901 8449 19935 8483
rect 22017 8449 22051 8483
rect 4537 8381 4571 8415
rect 7297 8381 7331 8415
rect 7757 8381 7791 8415
rect 9965 8381 9999 8415
rect 12449 8381 12483 8415
rect 15945 8381 15979 8415
rect 16773 8381 16807 8415
rect 17233 8381 17267 8415
rect 17509 8381 17543 8415
rect 23765 8381 23799 8415
rect 1685 8313 1719 8347
rect 2329 8313 2363 8347
rect 11713 8313 11747 8347
rect 15301 8313 15335 8347
rect 20637 8313 20671 8347
rect 21281 8313 21315 8347
rect 21833 8313 21867 8347
rect 25513 8313 25547 8347
rect 1961 8245 1995 8279
rect 3525 8245 3559 8279
rect 4813 8245 4847 8279
rect 4997 8245 5031 8279
rect 15025 8245 15059 8279
rect 18981 8245 19015 8279
rect 4261 8041 4295 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 9505 8041 9539 8075
rect 13737 8041 13771 8075
rect 16405 8041 16439 8075
rect 17969 8041 18003 8075
rect 18153 8041 18187 8075
rect 8493 7973 8527 8007
rect 8677 7973 8711 8007
rect 13461 7973 13495 8007
rect 17785 7973 17819 8007
rect 25329 7973 25363 8007
rect 1409 7905 1443 7939
rect 3893 7905 3927 7939
rect 7389 7905 7423 7939
rect 9045 7905 9079 7939
rect 13185 7905 13219 7939
rect 13645 7905 13679 7939
rect 14657 7905 14691 7939
rect 18705 7905 18739 7939
rect 21097 7905 21131 7939
rect 3985 7837 4019 7871
rect 4445 7837 4479 7871
rect 4537 7837 4571 7871
rect 6561 7837 6595 7871
rect 7021 7837 7055 7871
rect 8033 7837 8067 7871
rect 8585 7837 8619 7871
rect 9137 7837 9171 7871
rect 13921 7837 13955 7871
rect 20821 7837 20855 7871
rect 25053 7837 25087 7871
rect 25513 7837 25547 7871
rect 1685 7769 1719 7803
rect 6377 7769 6411 7803
rect 6837 7769 6871 7803
rect 14933 7769 14967 7803
rect 17509 7769 17543 7803
rect 18613 7769 18647 7803
rect 3157 7701 3191 7735
rect 6745 7701 6779 7735
rect 7205 7701 7239 7735
rect 18521 7701 18555 7735
rect 22569 7701 22603 7735
rect 25237 7701 25271 7735
rect 1593 7497 1627 7531
rect 2513 7497 2547 7531
rect 7297 7497 7331 7531
rect 11897 7497 11931 7531
rect 12817 7497 12851 7531
rect 15577 7497 15611 7531
rect 17325 7497 17359 7531
rect 1501 7429 1535 7463
rect 5917 7429 5951 7463
rect 6377 7429 6411 7463
rect 9505 7429 9539 7463
rect 9705 7429 9739 7463
rect 11989 7429 12023 7463
rect 15025 7429 15059 7463
rect 15853 7429 15887 7463
rect 22201 7429 22235 7463
rect 22293 7429 22327 7463
rect 25145 7429 25179 7463
rect 2605 7361 2639 7395
rect 6101 7361 6135 7395
rect 6193 7361 6227 7395
rect 6745 7361 6779 7395
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 8217 7361 8251 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9229 7361 9263 7395
rect 12357 7361 12391 7395
rect 12541 7361 12575 7395
rect 12633 7361 12667 7395
rect 15761 7361 15795 7395
rect 17417 7361 17451 7395
rect 17969 7361 18003 7395
rect 18521 7361 18555 7395
rect 18981 7361 19015 7395
rect 21373 7361 21407 7395
rect 2053 7293 2087 7327
rect 3065 7293 3099 7327
rect 6837 7293 6871 7327
rect 8493 7293 8527 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 12173 7293 12207 7327
rect 15485 7293 15519 7327
rect 16681 7293 16715 7327
rect 18245 7293 18279 7327
rect 22385 7293 22419 7327
rect 2421 7225 2455 7259
rect 2789 7225 2823 7259
rect 6193 7225 6227 7259
rect 7849 7225 7883 7259
rect 8309 7225 8343 7259
rect 9413 7225 9447 7259
rect 15393 7225 15427 7259
rect 16129 7225 16163 7259
rect 18153 7225 18187 7259
rect 21833 7225 21867 7259
rect 3709 7157 3743 7191
rect 7021 7157 7055 7191
rect 8953 7157 8987 7191
rect 9689 7157 9723 7191
rect 9873 7157 9907 7191
rect 11529 7157 11563 7191
rect 12633 7157 12667 7191
rect 16313 7157 16347 7191
rect 17509 7157 17543 7191
rect 17877 7157 17911 7191
rect 18061 7157 18095 7191
rect 18337 7157 18371 7191
rect 18797 7157 18831 7191
rect 21189 7157 21223 7191
rect 25421 7157 25455 7191
rect 7389 6953 7423 6987
rect 9229 6953 9263 6987
rect 10149 6953 10183 6987
rect 13185 6953 13219 6987
rect 18245 6953 18279 6987
rect 4169 6885 4203 6919
rect 4537 6885 4571 6919
rect 5089 6885 5123 6919
rect 9413 6885 9447 6919
rect 9873 6885 9907 6919
rect 11253 6885 11287 6919
rect 17969 6885 18003 6919
rect 18153 6885 18187 6919
rect 20269 6885 20303 6919
rect 5273 6817 5307 6851
rect 7665 6817 7699 6851
rect 9505 6817 9539 6851
rect 9965 6817 9999 6851
rect 18797 6817 18831 6851
rect 19349 6817 19383 6851
rect 22293 6817 22327 6851
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 5641 6749 5675 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 8585 6749 8619 6783
rect 8677 6749 8711 6783
rect 8953 6749 8987 6783
rect 10057 6749 10091 6783
rect 11437 6749 11471 6783
rect 16589 6749 16623 6783
rect 16773 6749 16807 6783
rect 17693 6749 17727 6783
rect 18613 6749 18647 6783
rect 20545 6749 20579 6783
rect 3893 6681 3927 6715
rect 4813 6681 4847 6715
rect 8309 6681 8343 6715
rect 10885 6681 10919 6715
rect 11713 6681 11747 6715
rect 19993 6681 20027 6715
rect 20821 6681 20855 6715
rect 4353 6613 4387 6647
rect 5457 6613 5491 6647
rect 6653 6613 6687 6647
rect 8033 6613 8067 6647
rect 10517 6613 10551 6647
rect 11345 6613 11379 6647
rect 16957 6613 16991 6647
rect 18705 6613 18739 6647
rect 19901 6613 19935 6647
rect 20453 6613 20487 6647
rect 7941 6409 7975 6443
rect 9137 6409 9171 6443
rect 11529 6409 11563 6443
rect 12357 6409 12391 6443
rect 14841 6409 14875 6443
rect 19809 6409 19843 6443
rect 20637 6409 20671 6443
rect 21465 6409 21499 6443
rect 8217 6341 8251 6375
rect 11805 6341 11839 6375
rect 15209 6341 15243 6375
rect 16681 6341 16715 6375
rect 18337 6341 18371 6375
rect 4537 6273 4571 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4905 6273 4939 6307
rect 5181 6273 5215 6307
rect 5641 6273 5675 6307
rect 5733 6273 5767 6307
rect 5825 6273 5859 6307
rect 6009 6273 6043 6307
rect 6837 6273 6871 6307
rect 7389 6273 7423 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8493 6273 8527 6307
rect 8585 6273 8619 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 9413 6273 9447 6307
rect 9597 6273 9631 6307
rect 9689 6273 9723 6307
rect 9873 6273 9907 6307
rect 10241 6273 10275 6307
rect 11713 6273 11747 6307
rect 12541 6273 12575 6307
rect 14381 6273 14415 6307
rect 15025 6273 15059 6307
rect 15301 6273 15335 6307
rect 15853 6273 15887 6307
rect 15946 6273 15980 6307
rect 16129 6273 16163 6307
rect 16221 6273 16255 6307
rect 16318 6273 16352 6307
rect 17601 6273 17635 6307
rect 20821 6273 20855 6307
rect 21649 6273 21683 6307
rect 22017 6273 22051 6307
rect 25237 6273 25271 6307
rect 7849 6205 7883 6239
rect 8769 6205 8803 6239
rect 9505 6205 9539 6239
rect 9965 6205 9999 6239
rect 10057 6205 10091 6239
rect 12265 6205 12299 6239
rect 14197 6205 14231 6239
rect 17509 6205 17543 6239
rect 18061 6205 18095 6239
rect 20913 6205 20947 6239
rect 21373 6205 21407 6239
rect 7297 6137 7331 6171
rect 12081 6137 12115 6171
rect 16497 6137 16531 6171
rect 17049 6137 17083 6171
rect 21189 6137 21223 6171
rect 25421 6137 25455 6171
rect 4261 6069 4295 6103
rect 4997 6069 5031 6103
rect 5365 6069 5399 6103
rect 6929 6069 6963 6103
rect 7573 6069 7607 6103
rect 10425 6069 10459 6103
rect 14565 6069 14599 6103
rect 17141 6069 17175 6103
rect 17877 6069 17911 6103
rect 21833 6069 21867 6103
rect 6653 5865 6687 5899
rect 7481 5865 7515 5899
rect 8585 5865 8619 5899
rect 15301 5865 15335 5899
rect 15393 5865 15427 5899
rect 17877 5865 17911 5899
rect 20821 5865 20855 5899
rect 7297 5797 7331 5831
rect 7849 5797 7883 5831
rect 8401 5797 8435 5831
rect 14565 5797 14599 5831
rect 14749 5797 14783 5831
rect 16865 5797 16899 5831
rect 19625 5797 19659 5831
rect 20637 5797 20671 5831
rect 5181 5729 5215 5763
rect 7021 5729 7055 5763
rect 7573 5729 7607 5763
rect 14657 5729 14691 5763
rect 15761 5729 15795 5763
rect 16405 5729 16439 5763
rect 19257 5729 19291 5763
rect 19717 5729 19751 5763
rect 20361 5729 20395 5763
rect 21189 5729 21223 5763
rect 4905 5661 4939 5695
rect 11805 5661 11839 5695
rect 13737 5661 13771 5695
rect 13921 5661 13955 5695
rect 14933 5661 14967 5695
rect 15025 5661 15059 5695
rect 15577 5661 15611 5695
rect 15669 5661 15703 5695
rect 15853 5661 15887 5695
rect 16483 5661 16517 5695
rect 17049 5661 17083 5695
rect 17233 5661 17267 5695
rect 17325 5661 17359 5695
rect 17785 5661 17819 5695
rect 18889 5661 18923 5695
rect 20913 5661 20947 5695
rect 1501 5593 1535 5627
rect 8125 5593 8159 5627
rect 14197 5593 14231 5627
rect 18521 5593 18555 5627
rect 18705 5593 18739 5627
rect 1593 5525 1627 5559
rect 8033 5525 8067 5559
rect 11621 5525 11655 5559
rect 13829 5525 13863 5559
rect 15117 5525 15151 5559
rect 16773 5525 16807 5559
rect 22661 5525 22695 5559
rect 7665 5321 7699 5355
rect 11161 5321 11195 5355
rect 16405 5321 16439 5355
rect 19533 5321 19567 5355
rect 20729 5321 20763 5355
rect 7849 5253 7883 5287
rect 11805 5253 11839 5287
rect 15393 5253 15427 5287
rect 16221 5253 16255 5287
rect 18245 5253 18279 5287
rect 20177 5253 20211 5287
rect 21833 5253 21867 5287
rect 1409 5185 1443 5219
rect 3985 5185 4019 5219
rect 7573 5185 7607 5219
rect 7757 5185 7791 5219
rect 11345 5185 11379 5219
rect 13829 5185 13863 5219
rect 13921 5185 13955 5219
rect 14013 5185 14047 5219
rect 14197 5185 14231 5219
rect 14657 5185 14691 5219
rect 15117 5185 15151 5219
rect 15209 5185 15243 5219
rect 15761 5185 15795 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 16497 5185 16531 5219
rect 21097 5185 21131 5219
rect 21189 5185 21223 5219
rect 25237 5185 25271 5219
rect 4261 5117 4295 5151
rect 11529 5117 11563 5151
rect 14749 5117 14783 5151
rect 15393 5117 15427 5151
rect 21373 5117 21407 5151
rect 20453 5049 20487 5083
rect 22109 5049 22143 5083
rect 1593 4981 1627 5015
rect 5733 4981 5767 5015
rect 9137 4981 9171 5015
rect 13277 4981 13311 5015
rect 13553 4981 13587 5015
rect 14933 4981 14967 5015
rect 15485 4981 15519 5015
rect 16221 4981 16255 5015
rect 20637 4981 20671 5015
rect 22293 4981 22327 5015
rect 25421 4981 25455 5015
rect 7573 4777 7607 4811
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 11253 4777 11287 4811
rect 14749 4777 14783 4811
rect 15485 4777 15519 4811
rect 15853 4777 15887 4811
rect 16037 4777 16071 4811
rect 16313 4777 16347 4811
rect 18705 4777 18739 4811
rect 8585 4709 8619 4743
rect 9873 4709 9907 4743
rect 13553 4709 13587 4743
rect 10057 4641 10091 4675
rect 11897 4641 11931 4675
rect 12633 4641 12667 4675
rect 13277 4641 13311 4675
rect 14105 4641 14139 4675
rect 1409 4573 1443 4607
rect 7481 4573 7515 4607
rect 8125 4573 8159 4607
rect 10333 4573 10367 4607
rect 11621 4573 11655 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 15301 4573 15335 4607
rect 15393 4573 15427 4607
rect 15945 4573 15979 4607
rect 16129 4573 16163 4607
rect 16221 4573 16255 4607
rect 16405 4573 16439 4607
rect 16957 4573 16991 4607
rect 21189 4573 21223 4607
rect 22017 4573 22051 4607
rect 25237 4573 25271 4607
rect 9597 4505 9631 4539
rect 17233 4505 17267 4539
rect 1593 4437 1627 4471
rect 10149 4437 10183 4471
rect 11713 4437 11747 4471
rect 13185 4437 13219 4471
rect 13737 4437 13771 4471
rect 14841 4437 14875 4471
rect 21005 4437 21039 4471
rect 22661 4437 22695 4471
rect 25421 4437 25455 4471
rect 14749 4233 14783 4267
rect 17877 4233 17911 4267
rect 5549 4097 5583 4131
rect 6377 4097 6411 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 8125 4097 8159 4131
rect 11069 4097 11103 4131
rect 13737 4097 13771 4131
rect 13921 4097 13955 4131
rect 14105 4097 14139 4131
rect 14657 4097 14691 4131
rect 14841 4097 14875 4131
rect 17325 4097 17359 4131
rect 18061 4097 18095 4131
rect 19901 4097 19935 4131
rect 22017 4097 22051 4131
rect 22293 4097 22327 4131
rect 7573 4029 7607 4063
rect 9045 4029 9079 4063
rect 9321 4029 9355 4063
rect 12541 4029 12575 4063
rect 13001 4029 13035 4063
rect 17785 4029 17819 4063
rect 20177 4029 20211 4063
rect 5917 3961 5951 3995
rect 6653 3961 6687 3995
rect 7849 3961 7883 3995
rect 10793 3961 10827 3995
rect 10885 3961 10919 3995
rect 12909 3961 12943 3995
rect 13737 3961 13771 3995
rect 14565 3961 14599 3995
rect 17601 3961 17635 3995
rect 21833 3961 21867 3995
rect 6009 3893 6043 3927
rect 6837 3893 6871 3927
rect 7021 3893 7055 3927
rect 7297 3893 7331 3927
rect 8033 3893 8067 3927
rect 8769 3893 8803 3927
rect 14197 3893 14231 3927
rect 21649 3893 21683 3927
rect 22109 3893 22143 3927
rect 2145 3689 2179 3723
rect 6364 3689 6398 3723
rect 7941 3689 7975 3723
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 11240 3689 11274 3723
rect 25053 3689 25087 3723
rect 7849 3621 7883 3655
rect 13185 3621 13219 3655
rect 13645 3621 13679 3655
rect 25329 3621 25363 3655
rect 6101 3553 6135 3587
rect 8401 3553 8435 3587
rect 8585 3553 8619 3587
rect 9597 3553 9631 3587
rect 10425 3553 10459 3587
rect 10977 3553 11011 3587
rect 21005 3553 21039 3587
rect 22753 3553 22787 3587
rect 22937 3553 22971 3587
rect 1961 3485 1995 3519
rect 4261 3485 4295 3519
rect 10149 3485 10183 3519
rect 10793 3485 10827 3519
rect 12817 3485 12851 3519
rect 13369 3485 13403 3519
rect 15117 3485 15151 3519
rect 15761 3485 15795 3519
rect 17785 3485 17819 3519
rect 20913 3485 20947 3519
rect 24777 3485 24811 3519
rect 25237 3485 25271 3519
rect 25513 3485 25547 3519
rect 1501 3417 1535 3451
rect 4537 3417 4571 3451
rect 8309 3417 8343 3451
rect 10241 3417 10275 3451
rect 16037 3417 16071 3451
rect 21281 3417 21315 3451
rect 1593 3349 1627 3383
rect 6009 3349 6043 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 10609 3349 10643 3383
rect 12725 3349 12759 3383
rect 13277 3349 13311 3383
rect 13829 3349 13863 3383
rect 14933 3349 14967 3383
rect 20729 3349 20763 3383
rect 23489 3349 23523 3383
rect 24961 3349 24995 3383
rect 5733 3145 5767 3179
rect 7205 3145 7239 3179
rect 15669 3145 15703 3179
rect 17233 3145 17267 3179
rect 20913 3145 20947 3179
rect 21833 3145 21867 3179
rect 22201 3145 22235 3179
rect 24409 3145 24443 3179
rect 1501 3077 1535 3111
rect 2605 3077 2639 3111
rect 11805 3077 11839 3111
rect 14197 3077 14231 3111
rect 16681 3077 16715 3111
rect 21373 3077 21407 3111
rect 22293 3077 22327 3111
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 3065 3009 3099 3043
rect 5917 3009 5951 3043
rect 6193 3009 6227 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 9873 3009 9907 3043
rect 10149 3009 10183 3043
rect 11529 3009 11563 3043
rect 13553 3009 13587 3043
rect 13921 3009 13955 3043
rect 17417 3009 17451 3043
rect 21281 3009 21315 3043
rect 24593 3009 24627 3043
rect 24777 3009 24811 3043
rect 25237 3009 25271 3043
rect 6837 2941 6871 2975
rect 7021 2941 7055 2975
rect 8309 2941 8343 2975
rect 9965 2941 9999 2975
rect 17141 2941 17175 2975
rect 21465 2941 21499 2975
rect 22385 2941 22419 2975
rect 3249 2873 3283 2907
rect 6009 2873 6043 2907
rect 6377 2873 6411 2907
rect 10333 2873 10367 2907
rect 13369 2873 13403 2907
rect 17049 2873 17083 2907
rect 1593 2805 1627 2839
rect 2697 2805 2731 2839
rect 9781 2805 9815 2839
rect 10149 2805 10183 2839
rect 13277 2805 13311 2839
rect 25053 2805 25087 2839
rect 25421 2805 25455 2839
rect 3157 2601 3191 2635
rect 4537 2601 4571 2635
rect 6561 2601 6595 2635
rect 9137 2601 9171 2635
rect 10609 2601 10643 2635
rect 12541 2601 12575 2635
rect 13645 2601 13679 2635
rect 15025 2601 15059 2635
rect 17233 2601 17267 2635
rect 21557 2601 21591 2635
rect 8033 2533 8067 2567
rect 14841 2533 14875 2567
rect 20269 2533 20303 2567
rect 24133 2533 24167 2567
rect 2145 2397 2179 2431
rect 2513 2397 2547 2431
rect 4353 2397 4387 2431
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 10425 2397 10459 2431
rect 11069 2397 11103 2431
rect 12265 2397 12299 2431
rect 12725 2397 12759 2431
rect 13093 2397 13127 2431
rect 13829 2397 13863 2431
rect 14565 2397 14599 2431
rect 15209 2397 15243 2431
rect 16773 2397 16807 2431
rect 17417 2397 17451 2431
rect 19809 2397 19843 2431
rect 20085 2397 20119 2431
rect 21281 2397 21315 2431
rect 21925 2397 21959 2431
rect 22661 2397 22695 2431
rect 22937 2397 22971 2431
rect 23949 2397 23983 2431
rect 25145 2397 25179 2431
rect 3065 2329 3099 2363
rect 3893 2329 3927 2363
rect 4721 2329 4755 2363
rect 5365 2329 5399 2363
rect 15761 2329 15795 2363
rect 18245 2329 18279 2363
rect 19349 2329 19383 2363
rect 24593 2329 24627 2363
rect 2605 2261 2639 2295
rect 4169 2261 4203 2295
rect 4813 2261 4847 2295
rect 5641 2261 5675 2295
rect 7389 2261 7423 2295
rect 9965 2261 9999 2295
rect 11253 2261 11287 2295
rect 12449 2261 12483 2295
rect 13185 2261 13219 2295
rect 15301 2261 15335 2295
rect 15853 2261 15887 2295
rect 16865 2261 16899 2295
rect 18337 2261 18371 2295
rect 19441 2261 19475 2295
rect 19993 2261 20027 2295
rect 22201 2261 22235 2295
rect 24869 2261 24903 2295
rect 25237 2261 25271 2295
<< metal1 >>
rect 1104 26682 25852 26704
rect 1104 26630 4043 26682
rect 4095 26630 4107 26682
rect 4159 26630 4171 26682
rect 4223 26630 4235 26682
rect 4287 26630 4299 26682
rect 4351 26630 10230 26682
rect 10282 26630 10294 26682
rect 10346 26630 10358 26682
rect 10410 26630 10422 26682
rect 10474 26630 10486 26682
rect 10538 26630 16417 26682
rect 16469 26630 16481 26682
rect 16533 26630 16545 26682
rect 16597 26630 16609 26682
rect 16661 26630 16673 26682
rect 16725 26630 22604 26682
rect 22656 26630 22668 26682
rect 22720 26630 22732 26682
rect 22784 26630 22796 26682
rect 22848 26630 22860 26682
rect 22912 26630 25852 26682
rect 1104 26608 25852 26630
rect 1578 26528 1584 26580
rect 1636 26528 1642 26580
rect 2222 26528 2228 26580
rect 2280 26528 2286 26580
rect 7374 26528 7380 26580
rect 7432 26528 7438 26580
rect 8386 26528 8392 26580
rect 8444 26568 8450 26580
rect 9125 26571 9183 26577
rect 9125 26568 9137 26571
rect 8444 26540 9137 26568
rect 8444 26528 8450 26540
rect 9125 26537 9137 26540
rect 9171 26537 9183 26571
rect 9125 26531 9183 26537
rect 11054 26528 11060 26580
rect 11112 26528 11118 26580
rect 11606 26528 11612 26580
rect 11664 26568 11670 26580
rect 11885 26571 11943 26577
rect 11885 26568 11897 26571
rect 11664 26540 11897 26568
rect 11664 26528 11670 26540
rect 11885 26537 11897 26540
rect 11931 26537 11943 26571
rect 11885 26531 11943 26537
rect 14458 26528 14464 26580
rect 14516 26528 14522 26580
rect 16758 26528 16764 26580
rect 16816 26568 16822 26580
rect 17037 26571 17095 26577
rect 17037 26568 17049 26571
rect 16816 26540 17049 26568
rect 16816 26528 16822 26540
rect 17037 26537 17049 26540
rect 17083 26537 17095 26571
rect 17678 26568 17684 26580
rect 17037 26531 17095 26537
rect 17420 26540 17684 26568
rect 3789 26503 3847 26509
rect 3789 26469 3801 26503
rect 3835 26500 3847 26503
rect 5902 26500 5908 26512
rect 3835 26472 5908 26500
rect 3835 26469 3847 26472
rect 3789 26463 3847 26469
rect 5902 26460 5908 26472
rect 5960 26460 5966 26512
rect 9953 26503 10011 26509
rect 9953 26469 9965 26503
rect 9999 26500 10011 26503
rect 10686 26500 10692 26512
rect 9999 26472 10692 26500
rect 9999 26469 10011 26472
rect 9953 26463 10011 26469
rect 10686 26460 10692 26472
rect 10744 26460 10750 26512
rect 15565 26503 15623 26509
rect 15565 26469 15577 26503
rect 15611 26500 15623 26503
rect 17420 26500 17448 26540
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 19058 26528 19064 26580
rect 19116 26568 19122 26580
rect 19429 26571 19487 26577
rect 19429 26568 19441 26571
rect 19116 26540 19441 26568
rect 19116 26528 19122 26540
rect 19429 26537 19441 26540
rect 19475 26537 19487 26571
rect 19429 26531 19487 26537
rect 19978 26528 19984 26580
rect 20036 26568 20042 26580
rect 20257 26571 20315 26577
rect 20257 26568 20269 26571
rect 20036 26540 20269 26568
rect 20036 26528 20042 26540
rect 20257 26537 20269 26540
rect 20303 26537 20315 26571
rect 20257 26531 20315 26537
rect 20714 26528 20720 26580
rect 20772 26568 20778 26580
rect 20901 26571 20959 26577
rect 20901 26568 20913 26571
rect 20772 26540 20913 26568
rect 20772 26528 20778 26540
rect 20901 26537 20913 26540
rect 20947 26537 20959 26571
rect 20901 26531 20959 26537
rect 23198 26528 23204 26580
rect 23256 26528 23262 26580
rect 23934 26528 23940 26580
rect 23992 26528 23998 26580
rect 15611 26472 17448 26500
rect 17497 26503 17555 26509
rect 15611 26469 15623 26472
rect 15565 26463 15623 26469
rect 17497 26469 17509 26503
rect 17543 26500 17555 26503
rect 18230 26500 18236 26512
rect 17543 26472 18236 26500
rect 17543 26469 17555 26472
rect 17497 26463 17555 26469
rect 18230 26460 18236 26472
rect 18288 26460 18294 26512
rect 18325 26503 18383 26509
rect 18325 26469 18337 26503
rect 18371 26469 18383 26503
rect 18325 26463 18383 26469
rect 22557 26503 22615 26509
rect 22557 26469 22569 26503
rect 22603 26500 22615 26503
rect 22830 26500 22836 26512
rect 22603 26472 22836 26500
rect 22603 26469 22615 26472
rect 22557 26463 22615 26469
rect 2682 26392 2688 26444
rect 2740 26392 2746 26444
rect 2884 26404 6868 26432
rect 1489 26299 1547 26305
rect 1489 26265 1501 26299
rect 1535 26296 1547 26299
rect 1762 26296 1768 26308
rect 1535 26268 1768 26296
rect 1535 26265 1547 26268
rect 1489 26259 1547 26265
rect 1762 26256 1768 26268
rect 1820 26256 1826 26308
rect 2133 26299 2191 26305
rect 2133 26265 2145 26299
rect 2179 26296 2191 26299
rect 2884 26296 2912 26404
rect 2961 26367 3019 26373
rect 2961 26333 2973 26367
rect 3007 26333 3019 26367
rect 2961 26327 3019 26333
rect 2179 26268 2912 26296
rect 2976 26296 3004 26327
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3292 26336 3985 26364
rect 3292 26324 3298 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 5166 26324 5172 26376
rect 5224 26364 5230 26376
rect 5261 26367 5319 26373
rect 5261 26364 5273 26367
rect 5224 26336 5273 26364
rect 5224 26324 5230 26336
rect 5261 26333 5273 26336
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5810 26324 5816 26376
rect 5868 26364 5874 26376
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5868 26336 5917 26364
rect 5868 26324 5874 26336
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6454 26324 6460 26376
rect 6512 26364 6518 26376
rect 6549 26367 6607 26373
rect 6549 26364 6561 26367
rect 6512 26336 6561 26364
rect 6512 26324 6518 26336
rect 6549 26333 6561 26336
rect 6595 26333 6607 26367
rect 6549 26327 6607 26333
rect 6840 26308 6868 26404
rect 17954 26392 17960 26444
rect 18012 26432 18018 26444
rect 18340 26432 18368 26463
rect 22830 26460 22836 26472
rect 22888 26460 22894 26512
rect 18012 26404 18368 26432
rect 23216 26432 23244 26528
rect 24854 26500 24860 26512
rect 23400 26472 24860 26500
rect 23216 26404 23336 26432
rect 18012 26392 18018 26404
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 9364 26336 9505 26364
rect 9364 26324 9370 26336
rect 9493 26333 9505 26336
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9674 26324 9680 26376
rect 9732 26364 9738 26376
rect 9769 26367 9827 26373
rect 9769 26364 9781 26367
rect 9732 26336 9781 26364
rect 9732 26324 9738 26336
rect 9769 26333 9781 26336
rect 9815 26333 9827 26367
rect 9769 26327 9827 26333
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12345 26367 12403 26373
rect 12345 26364 12357 26367
rect 12308 26336 12357 26364
rect 12308 26324 12314 26336
rect 12345 26333 12357 26336
rect 12391 26333 12403 26367
rect 12345 26327 12403 26333
rect 12894 26324 12900 26376
rect 12952 26364 12958 26376
rect 12989 26367 13047 26373
rect 12989 26364 13001 26367
rect 12952 26336 13001 26364
rect 12952 26324 12958 26336
rect 12989 26333 13001 26336
rect 13035 26333 13047 26367
rect 12989 26327 13047 26333
rect 15470 26324 15476 26376
rect 15528 26364 15534 26376
rect 15749 26367 15807 26373
rect 15749 26364 15761 26367
rect 15528 26336 15761 26364
rect 15528 26324 15534 26336
rect 15749 26333 15761 26336
rect 15795 26333 15807 26367
rect 16945 26367 17003 26373
rect 16945 26364 16957 26367
rect 15749 26327 15807 26333
rect 15856 26336 16957 26364
rect 3418 26296 3424 26308
rect 2976 26268 3424 26296
rect 2179 26265 2191 26268
rect 2133 26259 2191 26265
rect 3418 26256 3424 26268
rect 3476 26256 3482 26308
rect 6822 26256 6828 26308
rect 6880 26256 6886 26308
rect 7282 26256 7288 26308
rect 7340 26256 7346 26308
rect 8202 26256 8208 26308
rect 8260 26296 8266 26308
rect 9033 26299 9091 26305
rect 9033 26296 9045 26299
rect 8260 26268 9045 26296
rect 8260 26256 8266 26268
rect 9033 26265 9045 26268
rect 9079 26265 9091 26299
rect 9033 26259 9091 26265
rect 10226 26256 10232 26308
rect 10284 26296 10290 26308
rect 10965 26299 11023 26305
rect 10965 26296 10977 26299
rect 10284 26268 10977 26296
rect 10284 26256 10290 26268
rect 10965 26265 10977 26268
rect 11011 26265 11023 26299
rect 10965 26259 11023 26265
rect 11793 26299 11851 26305
rect 11793 26265 11805 26299
rect 11839 26296 11851 26299
rect 12066 26296 12072 26308
rect 11839 26268 12072 26296
rect 11839 26265 11851 26268
rect 11793 26259 11851 26265
rect 12066 26256 12072 26268
rect 12124 26256 12130 26308
rect 14090 26256 14096 26308
rect 14148 26296 14154 26308
rect 14369 26299 14427 26305
rect 14369 26296 14381 26299
rect 14148 26268 14381 26296
rect 14148 26256 14154 26268
rect 14369 26265 14381 26268
rect 14415 26265 14427 26299
rect 14369 26259 14427 26265
rect 15010 26256 15016 26308
rect 15068 26256 15074 26308
rect 15194 26256 15200 26308
rect 15252 26296 15258 26308
rect 15856 26296 15884 26336
rect 16945 26333 16957 26336
rect 16991 26333 17003 26367
rect 16945 26327 17003 26333
rect 17402 26324 17408 26376
rect 17460 26364 17466 26376
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 17460 26336 17693 26364
rect 17460 26324 17466 26336
rect 17681 26333 17693 26336
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 18046 26324 18052 26376
rect 18104 26364 18110 26376
rect 18141 26367 18199 26373
rect 18141 26364 18153 26367
rect 18104 26336 18153 26364
rect 18104 26324 18110 26336
rect 18141 26333 18153 26336
rect 18187 26333 18199 26367
rect 18141 26327 18199 26333
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 23308 26373 23336 26404
rect 22373 26367 22431 26373
rect 22373 26364 22385 26367
rect 22152 26336 22385 26364
rect 22152 26324 22158 26336
rect 22373 26333 22385 26336
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 23201 26367 23259 26373
rect 23201 26333 23213 26367
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26333 23351 26367
rect 23293 26327 23351 26333
rect 15252 26268 15884 26296
rect 15252 26256 15258 26268
rect 16850 26256 16856 26308
rect 16908 26296 16914 26308
rect 19337 26299 19395 26305
rect 19337 26296 19349 26299
rect 16908 26268 19349 26296
rect 16908 26256 16914 26268
rect 19337 26265 19349 26268
rect 19383 26265 19395 26299
rect 19337 26259 19395 26265
rect 19426 26256 19432 26308
rect 19484 26296 19490 26308
rect 20165 26299 20223 26305
rect 20165 26296 20177 26299
rect 19484 26268 20177 26296
rect 19484 26256 19490 26268
rect 20165 26265 20177 26268
rect 20211 26265 20223 26299
rect 20165 26259 20223 26265
rect 20809 26299 20867 26305
rect 20809 26265 20821 26299
rect 20855 26296 20867 26299
rect 21726 26296 21732 26308
rect 20855 26268 21732 26296
rect 20855 26265 20867 26268
rect 20809 26259 20867 26265
rect 21726 26256 21732 26268
rect 21784 26256 21790 26308
rect 21910 26256 21916 26308
rect 21968 26256 21974 26308
rect 23216 26296 23244 26327
rect 23400 26296 23428 26472
rect 24854 26460 24860 26472
rect 24912 26460 24918 26512
rect 24578 26392 24584 26444
rect 24636 26392 24642 26444
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 25866 26364 25872 26376
rect 24903 26336 25872 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 25866 26324 25872 26336
rect 25924 26324 25930 26376
rect 23216 26268 23428 26296
rect 23842 26256 23848 26308
rect 23900 26256 23906 26308
rect 5442 26188 5448 26240
rect 5500 26188 5506 26240
rect 6086 26188 6092 26240
rect 6144 26188 6150 26240
rect 6730 26188 6736 26240
rect 6788 26188 6794 26240
rect 9674 26188 9680 26240
rect 9732 26188 9738 26240
rect 12529 26231 12587 26237
rect 12529 26197 12541 26231
rect 12575 26228 12587 26231
rect 12618 26228 12624 26240
rect 12575 26200 12624 26228
rect 12575 26197 12587 26200
rect 12529 26191 12587 26197
rect 12618 26188 12624 26200
rect 12676 26188 12682 26240
rect 13170 26188 13176 26240
rect 13228 26188 13234 26240
rect 14826 26188 14832 26240
rect 14884 26228 14890 26240
rect 15105 26231 15163 26237
rect 15105 26228 15117 26231
rect 14884 26200 15117 26228
rect 14884 26188 14890 26200
rect 15105 26197 15117 26200
rect 15151 26197 15163 26231
rect 15105 26191 15163 26197
rect 21266 26188 21272 26240
rect 21324 26228 21330 26240
rect 22005 26231 22063 26237
rect 22005 26228 22017 26231
rect 21324 26200 22017 26228
rect 21324 26188 21330 26200
rect 22005 26197 22017 26200
rect 22051 26197 22063 26231
rect 22005 26191 22063 26197
rect 23014 26188 23020 26240
rect 23072 26188 23078 26240
rect 23106 26188 23112 26240
rect 23164 26228 23170 26240
rect 23477 26231 23535 26237
rect 23477 26228 23489 26231
rect 23164 26200 23489 26228
rect 23164 26188 23170 26200
rect 23477 26197 23489 26200
rect 23523 26197 23535 26231
rect 23477 26191 23535 26197
rect 1104 26138 25852 26160
rect 1104 26086 4703 26138
rect 4755 26086 4767 26138
rect 4819 26086 4831 26138
rect 4883 26086 4895 26138
rect 4947 26086 4959 26138
rect 5011 26086 10890 26138
rect 10942 26086 10954 26138
rect 11006 26086 11018 26138
rect 11070 26086 11082 26138
rect 11134 26086 11146 26138
rect 11198 26086 17077 26138
rect 17129 26086 17141 26138
rect 17193 26086 17205 26138
rect 17257 26086 17269 26138
rect 17321 26086 17333 26138
rect 17385 26086 23264 26138
rect 23316 26086 23328 26138
rect 23380 26086 23392 26138
rect 23444 26086 23456 26138
rect 23508 26086 23520 26138
rect 23572 26086 25852 26138
rect 1104 26064 25852 26086
rect 1026 25984 1032 26036
rect 1084 26024 1090 26036
rect 1949 26027 2007 26033
rect 1949 26024 1961 26027
rect 1084 25996 1961 26024
rect 1084 25984 1090 25996
rect 1949 25993 1961 25996
rect 1995 25993 2007 26027
rect 1949 25987 2007 25993
rect 5902 25984 5908 26036
rect 5960 26024 5966 26036
rect 7837 26027 7895 26033
rect 7837 26024 7849 26027
rect 5960 25996 7849 26024
rect 5960 25984 5966 25996
rect 7837 25993 7849 25996
rect 7883 25993 7895 26027
rect 7837 25987 7895 25993
rect 7929 26027 7987 26033
rect 7929 25993 7941 26027
rect 7975 26024 7987 26027
rect 7975 25996 12434 26024
rect 7975 25993 7987 25996
rect 7929 25987 7987 25993
rect 658 25916 664 25968
rect 716 25956 722 25968
rect 8570 25956 8576 25968
rect 716 25928 3188 25956
rect 716 25916 722 25928
rect 1854 25848 1860 25900
rect 1912 25848 1918 25900
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25857 2467 25891
rect 2409 25851 2467 25857
rect 2424 25752 2452 25851
rect 2866 25848 2872 25900
rect 2924 25848 2930 25900
rect 3160 25897 3188 25928
rect 7484 25928 8576 25956
rect 3145 25891 3203 25897
rect 3145 25857 3157 25891
rect 3191 25857 3203 25891
rect 3145 25851 3203 25857
rect 7484 25752 7512 25928
rect 8570 25916 8576 25928
rect 8628 25916 8634 25968
rect 9030 25916 9036 25968
rect 9088 25916 9094 25968
rect 10134 25916 10140 25968
rect 10192 25956 10198 25968
rect 10192 25928 11744 25956
rect 10192 25916 10198 25928
rect 10226 25848 10232 25900
rect 10284 25848 10290 25900
rect 11716 25897 11744 25928
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11974 25848 11980 25900
rect 12032 25848 12038 25900
rect 8110 25780 8116 25832
rect 8168 25780 8174 25832
rect 8294 25780 8300 25832
rect 8352 25780 8358 25832
rect 8573 25823 8631 25829
rect 8573 25789 8585 25823
rect 8619 25820 8631 25823
rect 8662 25820 8668 25832
rect 8619 25792 8668 25820
rect 8619 25789 8631 25792
rect 8573 25783 8631 25789
rect 8662 25780 8668 25792
rect 8720 25780 8726 25832
rect 10045 25823 10103 25829
rect 10045 25789 10057 25823
rect 10091 25820 10103 25823
rect 10244 25820 10272 25848
rect 10091 25792 10272 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10870 25780 10876 25832
rect 10928 25780 10934 25832
rect 11241 25755 11299 25761
rect 2424 25724 7512 25752
rect 9600 25724 10916 25752
rect 14 25644 20 25696
rect 72 25684 78 25696
rect 2501 25687 2559 25693
rect 2501 25684 2513 25687
rect 72 25656 2513 25684
rect 72 25644 78 25656
rect 2501 25653 2513 25656
rect 2547 25653 2559 25687
rect 2501 25647 2559 25653
rect 3050 25644 3056 25696
rect 3108 25644 3114 25696
rect 3326 25644 3332 25696
rect 3384 25644 3390 25696
rect 7469 25687 7527 25693
rect 7469 25653 7481 25687
rect 7515 25684 7527 25687
rect 8570 25684 8576 25696
rect 7515 25656 8576 25684
rect 7515 25653 7527 25656
rect 7469 25647 7527 25653
rect 8570 25644 8576 25656
rect 8628 25644 8634 25696
rect 8938 25644 8944 25696
rect 8996 25684 9002 25696
rect 9600 25684 9628 25724
rect 8996 25656 9628 25684
rect 8996 25644 9002 25656
rect 10594 25644 10600 25696
rect 10652 25684 10658 25696
rect 10781 25687 10839 25693
rect 10781 25684 10793 25687
rect 10652 25656 10793 25684
rect 10652 25644 10658 25656
rect 10781 25653 10793 25656
rect 10827 25653 10839 25687
rect 10888 25684 10916 25724
rect 11241 25721 11253 25755
rect 11287 25752 11299 25755
rect 11422 25752 11428 25764
rect 11287 25724 11428 25752
rect 11287 25721 11299 25724
rect 11241 25715 11299 25721
rect 11422 25712 11428 25724
rect 11480 25712 11486 25764
rect 12406 25752 12434 25996
rect 16206 25984 16212 26036
rect 16264 26024 16270 26036
rect 16301 26027 16359 26033
rect 16301 26024 16313 26027
rect 16264 25996 16313 26024
rect 16264 25984 16270 25996
rect 16301 25993 16313 25996
rect 16347 25993 16359 26027
rect 16301 25987 16359 25993
rect 17589 26027 17647 26033
rect 17589 25993 17601 26027
rect 17635 26024 17647 26027
rect 20993 26027 21051 26033
rect 17635 25996 18184 26024
rect 17635 25993 17647 25996
rect 17589 25987 17647 25993
rect 18156 25965 18184 25996
rect 20993 25993 21005 26027
rect 21039 26024 21051 26027
rect 23014 26024 23020 26036
rect 21039 25996 23020 26024
rect 21039 25993 21051 25996
rect 20993 25987 21051 25993
rect 23014 25984 23020 25996
rect 23072 25984 23078 26036
rect 18141 25959 18199 25965
rect 18141 25925 18153 25959
rect 18187 25925 18199 25959
rect 18141 25919 18199 25925
rect 18782 25916 18788 25968
rect 18840 25916 18846 25968
rect 24213 25959 24271 25965
rect 24213 25956 24225 25959
rect 19628 25928 24225 25956
rect 15930 25848 15936 25900
rect 15988 25888 15994 25900
rect 16209 25891 16267 25897
rect 16209 25888 16221 25891
rect 15988 25860 16221 25888
rect 15988 25848 15994 25860
rect 16209 25857 16221 25860
rect 16255 25857 16267 25891
rect 16209 25851 16267 25857
rect 16393 25891 16451 25897
rect 16393 25857 16405 25891
rect 16439 25857 16451 25891
rect 16393 25851 16451 25857
rect 16114 25780 16120 25832
rect 16172 25820 16178 25832
rect 16408 25820 16436 25851
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 16172 25792 16436 25820
rect 16172 25780 16178 25792
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 19628 25829 19656 25928
rect 24213 25925 24225 25928
rect 24259 25925 24271 25959
rect 24213 25919 24271 25925
rect 20346 25848 20352 25900
rect 20404 25888 20410 25900
rect 21637 25891 21695 25897
rect 21637 25888 21649 25891
rect 20404 25860 21649 25888
rect 20404 25848 20410 25860
rect 21637 25857 21649 25860
rect 21683 25857 21695 25891
rect 21637 25851 21695 25857
rect 22922 25848 22928 25900
rect 22980 25888 22986 25900
rect 23753 25891 23811 25897
rect 23753 25888 23765 25891
rect 22980 25860 23765 25888
rect 22980 25848 22986 25860
rect 23753 25857 23765 25860
rect 23799 25857 23811 25891
rect 23753 25851 23811 25857
rect 24581 25891 24639 25897
rect 24581 25857 24593 25891
rect 24627 25888 24639 25891
rect 25314 25888 25320 25900
rect 24627 25860 25320 25888
rect 24627 25857 24639 25860
rect 24581 25851 24639 25857
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 26418 25848 26424 25900
rect 26476 25848 26482 25900
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 17972 25792 19625 25820
rect 17972 25752 18000 25792
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 19702 25780 19708 25832
rect 19760 25820 19766 25832
rect 21085 25823 21143 25829
rect 21085 25820 21097 25823
rect 19760 25792 21097 25820
rect 19760 25780 19766 25792
rect 21085 25789 21097 25792
rect 21131 25789 21143 25823
rect 21085 25783 21143 25789
rect 21177 25823 21235 25829
rect 21177 25789 21189 25823
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 24673 25823 24731 25829
rect 24673 25789 24685 25823
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 21192 25752 21220 25783
rect 21542 25752 21548 25764
rect 12406 25724 18000 25752
rect 20548 25724 21548 25752
rect 11333 25687 11391 25693
rect 11333 25684 11345 25687
rect 10888 25656 11345 25684
rect 10781 25647 10839 25653
rect 11333 25653 11345 25656
rect 11379 25653 11391 25687
rect 11333 25647 11391 25653
rect 11514 25644 11520 25696
rect 11572 25644 11578 25696
rect 11790 25644 11796 25696
rect 11848 25644 11854 25696
rect 18506 25644 18512 25696
rect 18564 25684 18570 25696
rect 20548 25684 20576 25724
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 24688 25752 24716 25783
rect 24946 25780 24952 25832
rect 25004 25780 25010 25832
rect 26436 25752 26464 25848
rect 24688 25724 26464 25752
rect 18564 25656 20576 25684
rect 20625 25687 20683 25693
rect 18564 25644 18570 25656
rect 20625 25653 20637 25687
rect 20671 25684 20683 25687
rect 21174 25684 21180 25696
rect 20671 25656 21180 25684
rect 20671 25653 20683 25656
rect 20625 25647 20683 25653
rect 21174 25644 21180 25656
rect 21232 25644 21238 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 23934 25644 23940 25696
rect 23992 25644 23998 25696
rect 1104 25594 25852 25616
rect 1104 25542 4043 25594
rect 4095 25542 4107 25594
rect 4159 25542 4171 25594
rect 4223 25542 4235 25594
rect 4287 25542 4299 25594
rect 4351 25542 10230 25594
rect 10282 25542 10294 25594
rect 10346 25542 10358 25594
rect 10410 25542 10422 25594
rect 10474 25542 10486 25594
rect 10538 25542 16417 25594
rect 16469 25542 16481 25594
rect 16533 25542 16545 25594
rect 16597 25542 16609 25594
rect 16661 25542 16673 25594
rect 16725 25542 22604 25594
rect 22656 25542 22668 25594
rect 22720 25542 22732 25594
rect 22784 25542 22796 25594
rect 22848 25542 22860 25594
rect 22912 25542 25852 25594
rect 1104 25520 25852 25542
rect 1394 25440 1400 25492
rect 1452 25480 1458 25492
rect 1581 25483 1639 25489
rect 1581 25480 1593 25483
rect 1452 25452 1593 25480
rect 1452 25440 1458 25452
rect 1581 25449 1593 25452
rect 1627 25449 1639 25483
rect 1581 25443 1639 25449
rect 8202 25440 8208 25492
rect 8260 25440 8266 25492
rect 8941 25483 8999 25489
rect 8941 25449 8953 25483
rect 8987 25480 8999 25483
rect 9030 25480 9036 25492
rect 8987 25452 9036 25480
rect 8987 25449 8999 25452
rect 8941 25443 8999 25449
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 9769 25483 9827 25489
rect 9769 25449 9781 25483
rect 9815 25480 9827 25483
rect 10134 25480 10140 25492
rect 9815 25452 10140 25480
rect 9815 25449 9827 25452
rect 9769 25443 9827 25449
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 11422 25480 11428 25492
rect 10888 25452 11428 25480
rect 8110 25372 8116 25424
rect 8168 25412 8174 25424
rect 9585 25415 9643 25421
rect 8168 25384 9536 25412
rect 8168 25372 8174 25384
rect 6457 25347 6515 25353
rect 6457 25313 6469 25347
rect 6503 25344 6515 25347
rect 8294 25344 8300 25356
rect 6503 25316 8300 25344
rect 6503 25313 6515 25316
rect 6457 25307 6515 25313
rect 8294 25304 8300 25316
rect 8352 25344 8358 25356
rect 9508 25344 9536 25384
rect 9585 25381 9597 25415
rect 9631 25412 9643 25415
rect 10888 25412 10916 25452
rect 11422 25440 11428 25452
rect 11480 25440 11486 25492
rect 12529 25483 12587 25489
rect 12529 25449 12541 25483
rect 12575 25480 12587 25483
rect 12894 25480 12900 25492
rect 12575 25452 12900 25480
rect 12575 25449 12587 25452
rect 12529 25443 12587 25449
rect 12894 25440 12900 25452
rect 12952 25480 12958 25492
rect 12952 25452 15516 25480
rect 12952 25440 12958 25452
rect 9631 25384 10916 25412
rect 9631 25381 9643 25384
rect 9585 25375 9643 25381
rect 12802 25372 12808 25424
rect 12860 25412 12866 25424
rect 12989 25415 13047 25421
rect 12989 25412 13001 25415
rect 12860 25384 13001 25412
rect 12860 25372 12866 25384
rect 12989 25381 13001 25384
rect 13035 25381 13047 25415
rect 12989 25375 13047 25381
rect 13173 25415 13231 25421
rect 13173 25381 13185 25415
rect 13219 25412 13231 25415
rect 13814 25412 13820 25424
rect 13219 25384 13820 25412
rect 13219 25381 13231 25384
rect 13173 25375 13231 25381
rect 13814 25372 13820 25384
rect 13872 25372 13878 25424
rect 15488 25412 15516 25452
rect 15838 25440 15844 25492
rect 15896 25440 15902 25492
rect 16850 25440 16856 25492
rect 16908 25440 16914 25492
rect 17402 25440 17408 25492
rect 17460 25440 17466 25492
rect 17770 25440 17776 25492
rect 17828 25480 17834 25492
rect 17865 25483 17923 25489
rect 17865 25480 17877 25483
rect 17828 25452 17877 25480
rect 17828 25440 17834 25452
rect 17865 25449 17877 25452
rect 17911 25449 17923 25483
rect 17865 25443 17923 25449
rect 18782 25440 18788 25492
rect 18840 25440 18846 25492
rect 19702 25480 19708 25492
rect 18892 25452 19708 25480
rect 18892 25412 18920 25452
rect 19702 25440 19708 25452
rect 19760 25440 19766 25492
rect 20346 25440 20352 25492
rect 20404 25440 20410 25492
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 25409 25483 25467 25489
rect 25409 25449 25421 25483
rect 25455 25480 25467 25483
rect 25498 25480 25504 25492
rect 25455 25452 25504 25480
rect 25455 25449 25467 25452
rect 25409 25443 25467 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 15488 25384 18920 25412
rect 19613 25415 19671 25421
rect 19613 25381 19625 25415
rect 19659 25412 19671 25415
rect 20070 25412 20076 25424
rect 19659 25384 20076 25412
rect 19659 25381 19671 25384
rect 19613 25375 19671 25381
rect 20070 25372 20076 25384
rect 20128 25412 20134 25424
rect 20165 25415 20223 25421
rect 20165 25412 20177 25415
rect 20128 25384 20177 25412
rect 20128 25372 20134 25384
rect 20165 25381 20177 25384
rect 20211 25381 20223 25415
rect 20165 25375 20223 25381
rect 10410 25344 10416 25356
rect 8352 25316 9444 25344
rect 9508 25316 10416 25344
rect 8352 25304 8358 25316
rect 1026 25236 1032 25288
rect 1084 25276 1090 25288
rect 1949 25279 2007 25285
rect 1949 25276 1961 25279
rect 1084 25248 1961 25276
rect 1084 25236 1090 25248
rect 1949 25245 1961 25248
rect 1995 25245 2007 25279
rect 1949 25239 2007 25245
rect 6362 25236 6368 25288
rect 6420 25236 6426 25288
rect 8481 25279 8539 25285
rect 8481 25245 8493 25279
rect 8527 25245 8539 25279
rect 8481 25239 8539 25245
rect 1489 25211 1547 25217
rect 1489 25177 1501 25211
rect 1535 25208 1547 25211
rect 2038 25208 2044 25220
rect 1535 25180 2044 25208
rect 1535 25177 1547 25180
rect 1489 25171 1547 25177
rect 2038 25168 2044 25180
rect 2096 25168 2102 25220
rect 6733 25211 6791 25217
rect 6733 25208 6745 25211
rect 6196 25180 6745 25208
rect 2133 25143 2191 25149
rect 2133 25109 2145 25143
rect 2179 25140 2191 25143
rect 2682 25140 2688 25152
rect 2179 25112 2688 25140
rect 2179 25109 2191 25112
rect 2133 25103 2191 25109
rect 2682 25100 2688 25112
rect 2740 25100 2746 25152
rect 6196 25149 6224 25180
rect 6733 25177 6745 25180
rect 6779 25177 6791 25211
rect 8496 25208 8524 25239
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 8757 25279 8815 25285
rect 8757 25276 8769 25279
rect 8628 25248 8769 25276
rect 8628 25236 8634 25248
rect 8757 25245 8769 25248
rect 8803 25245 8815 25279
rect 8757 25239 8815 25245
rect 8938 25236 8944 25288
rect 8996 25236 9002 25288
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9416 25276 9444 25316
rect 10410 25304 10416 25316
rect 10468 25304 10474 25356
rect 11057 25347 11115 25353
rect 11057 25313 11069 25347
rect 11103 25344 11115 25347
rect 11514 25344 11520 25356
rect 11103 25316 11520 25344
rect 11103 25313 11115 25316
rect 11057 25307 11115 25313
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 13722 25304 13728 25356
rect 13780 25344 13786 25356
rect 14093 25347 14151 25353
rect 14093 25344 14105 25347
rect 13780 25316 14105 25344
rect 13780 25304 13786 25316
rect 14093 25313 14105 25316
rect 14139 25344 14151 25347
rect 17862 25344 17868 25356
rect 14139 25316 17868 25344
rect 14139 25313 14151 25316
rect 14093 25307 14151 25313
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 18506 25304 18512 25356
rect 18564 25304 18570 25356
rect 19705 25347 19763 25353
rect 19705 25344 19717 25347
rect 18984 25316 19717 25344
rect 10781 25279 10839 25285
rect 9416 25272 10732 25276
rect 10781 25272 10793 25279
rect 9416 25248 10793 25272
rect 9125 25239 9183 25245
rect 8956 25208 8984 25236
rect 7958 25180 8340 25208
rect 8496 25180 8984 25208
rect 6733 25171 6791 25177
rect 8312 25149 8340 25180
rect 6181 25143 6239 25149
rect 6181 25109 6193 25143
rect 6227 25109 6239 25143
rect 6181 25103 6239 25109
rect 8297 25143 8355 25149
rect 8297 25109 8309 25143
rect 8343 25109 8355 25143
rect 8297 25103 8355 25109
rect 8570 25100 8576 25152
rect 8628 25100 8634 25152
rect 9140 25140 9168 25239
rect 9217 25211 9275 25217
rect 9217 25177 9229 25211
rect 9263 25208 9275 25211
rect 9766 25208 9772 25220
rect 9263 25180 9772 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 10229 25211 10287 25217
rect 10229 25177 10241 25211
rect 10275 25208 10287 25211
rect 10502 25208 10508 25220
rect 10275 25180 10508 25208
rect 10275 25177 10287 25180
rect 10229 25171 10287 25177
rect 10502 25168 10508 25180
rect 10560 25168 10566 25220
rect 9677 25143 9735 25149
rect 9677 25140 9689 25143
rect 9140 25112 9689 25140
rect 9677 25109 9689 25112
rect 9723 25109 9735 25143
rect 9677 25103 9735 25109
rect 10134 25100 10140 25152
rect 10192 25100 10198 25152
rect 10612 25140 10640 25248
rect 10704 25245 10793 25248
rect 10827 25245 10839 25279
rect 10704 25244 10839 25245
rect 10781 25239 10839 25244
rect 13170 25236 13176 25288
rect 13228 25276 13234 25288
rect 13909 25279 13967 25285
rect 13909 25276 13921 25279
rect 13228 25248 13921 25276
rect 13228 25236 13234 25248
rect 13909 25245 13921 25248
rect 13955 25245 13967 25279
rect 13909 25239 13967 25245
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16666 25276 16672 25288
rect 16163 25248 16672 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 11790 25168 11796 25220
rect 11848 25168 11854 25220
rect 12710 25168 12716 25220
rect 12768 25168 12774 25220
rect 14366 25168 14372 25220
rect 14424 25168 14430 25220
rect 16132 25208 16160 25239
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17313 25279 17371 25285
rect 17313 25276 17325 25279
rect 16807 25248 16896 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 14476 25180 14858 25208
rect 15672 25180 16160 25208
rect 11238 25140 11244 25152
rect 10612 25112 11244 25140
rect 11238 25100 11244 25112
rect 11296 25100 11302 25152
rect 13725 25143 13783 25149
rect 13725 25109 13737 25143
rect 13771 25140 13783 25143
rect 14476 25140 14504 25180
rect 13771 25112 14504 25140
rect 13771 25109 13783 25112
rect 13725 25103 13783 25109
rect 15102 25100 15108 25152
rect 15160 25140 15166 25152
rect 15672 25140 15700 25180
rect 16868 25152 16896 25248
rect 17236 25248 17325 25276
rect 15160 25112 15700 25140
rect 15160 25100 15166 25112
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 16669 25143 16727 25149
rect 16669 25140 16681 25143
rect 16632 25112 16681 25140
rect 16632 25100 16638 25112
rect 16669 25109 16681 25112
rect 16715 25109 16727 25143
rect 16669 25103 16727 25109
rect 16850 25100 16856 25152
rect 16908 25100 16914 25152
rect 16942 25100 16948 25152
rect 17000 25140 17006 25152
rect 17236 25149 17264 25248
rect 17313 25245 17325 25248
rect 17359 25245 17371 25279
rect 17313 25239 17371 25245
rect 18230 25236 18236 25288
rect 18288 25236 18294 25288
rect 18984 25285 19012 25316
rect 19705 25313 19717 25316
rect 19751 25313 19763 25347
rect 25774 25344 25780 25356
rect 19705 25307 19763 25313
rect 24228 25316 25780 25344
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25245 19027 25279
rect 18969 25239 19027 25245
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 24228 25285 24256 25316
rect 25774 25304 25780 25316
rect 25832 25304 25838 25356
rect 20441 25279 20499 25285
rect 20441 25276 20453 25279
rect 19392 25248 20453 25276
rect 19392 25236 19398 25248
rect 20441 25245 20453 25248
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 24213 25279 24271 25285
rect 24213 25245 24225 25279
rect 24259 25245 24271 25279
rect 24213 25239 24271 25245
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24544 25248 24685 25276
rect 24544 25236 24550 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 19245 25211 19303 25217
rect 19245 25177 19257 25211
rect 19291 25208 19303 25211
rect 19518 25208 19524 25220
rect 19291 25180 19524 25208
rect 19291 25177 19303 25180
rect 19245 25171 19303 25177
rect 19518 25168 19524 25180
rect 19576 25208 19582 25220
rect 19889 25211 19947 25217
rect 19889 25208 19901 25211
rect 19576 25180 19901 25208
rect 19576 25168 19582 25180
rect 19889 25177 19901 25180
rect 19935 25177 19947 25211
rect 20717 25211 20775 25217
rect 19889 25171 19947 25177
rect 20272 25180 20484 25208
rect 17221 25143 17279 25149
rect 17221 25140 17233 25143
rect 17000 25112 17233 25140
rect 17000 25100 17006 25112
rect 17221 25109 17233 25112
rect 17267 25109 17279 25143
rect 17221 25103 17279 25109
rect 17770 25100 17776 25152
rect 17828 25100 17834 25152
rect 18325 25143 18383 25149
rect 18325 25109 18337 25143
rect 18371 25140 18383 25143
rect 20272 25140 20300 25180
rect 18371 25112 20300 25140
rect 20456 25140 20484 25180
rect 20717 25177 20729 25211
rect 20763 25208 20775 25211
rect 20990 25208 20996 25220
rect 20763 25180 20996 25208
rect 20763 25177 20775 25180
rect 20717 25171 20775 25177
rect 20990 25168 20996 25180
rect 21048 25168 21054 25220
rect 21450 25168 21456 25220
rect 21508 25168 21514 25220
rect 25133 25211 25191 25217
rect 22112 25180 23796 25208
rect 22112 25140 22140 25180
rect 23768 25152 23796 25180
rect 25133 25177 25145 25211
rect 25179 25208 25191 25211
rect 26142 25208 26148 25220
rect 25179 25180 26148 25208
rect 25179 25177 25191 25180
rect 25133 25171 25191 25177
rect 26142 25168 26148 25180
rect 26200 25168 26206 25220
rect 20456 25112 22140 25140
rect 18371 25109 18383 25112
rect 18325 25103 18383 25109
rect 22186 25100 22192 25152
rect 22244 25100 22250 25152
rect 23750 25100 23756 25152
rect 23808 25100 23814 25152
rect 24026 25100 24032 25152
rect 24084 25100 24090 25152
rect 1104 25050 25852 25072
rect 1104 24998 4703 25050
rect 4755 24998 4767 25050
rect 4819 24998 4831 25050
rect 4883 24998 4895 25050
rect 4947 24998 4959 25050
rect 5011 24998 10890 25050
rect 10942 24998 10954 25050
rect 11006 24998 11018 25050
rect 11070 24998 11082 25050
rect 11134 24998 11146 25050
rect 11198 24998 17077 25050
rect 17129 24998 17141 25050
rect 17193 24998 17205 25050
rect 17257 24998 17269 25050
rect 17321 24998 17333 25050
rect 17385 24998 23264 25050
rect 23316 24998 23328 25050
rect 23380 24998 23392 25050
rect 23444 24998 23456 25050
rect 23508 24998 23520 25050
rect 23572 24998 25852 25050
rect 1104 24976 25852 24998
rect 6362 24896 6368 24948
rect 6420 24896 6426 24948
rect 11974 24896 11980 24948
rect 12032 24896 12038 24948
rect 13170 24896 13176 24948
rect 13228 24896 13234 24948
rect 14366 24896 14372 24948
rect 14424 24936 14430 24948
rect 15105 24939 15163 24945
rect 15105 24936 15117 24939
rect 14424 24908 15117 24936
rect 14424 24896 14430 24908
rect 15105 24905 15117 24908
rect 15151 24905 15163 24939
rect 15105 24899 15163 24905
rect 15286 24896 15292 24948
rect 15344 24936 15350 24948
rect 16393 24939 16451 24945
rect 16393 24936 16405 24939
rect 15344 24908 16405 24936
rect 15344 24896 15350 24908
rect 16393 24905 16405 24908
rect 16439 24905 16451 24939
rect 16393 24899 16451 24905
rect 16574 24896 16580 24948
rect 16632 24896 16638 24948
rect 17129 24939 17187 24945
rect 17129 24905 17141 24939
rect 17175 24936 17187 24939
rect 17402 24936 17408 24948
rect 17175 24908 17408 24936
rect 17175 24905 17187 24908
rect 17129 24899 17187 24905
rect 17402 24896 17408 24908
rect 17460 24896 17466 24948
rect 19426 24896 19432 24948
rect 19484 24896 19490 24948
rect 20990 24896 20996 24948
rect 21048 24936 21054 24948
rect 21453 24939 21511 24945
rect 21453 24936 21465 24939
rect 21048 24908 21465 24936
rect 21048 24896 21054 24908
rect 21453 24905 21465 24908
rect 21499 24905 21511 24939
rect 21453 24899 21511 24905
rect 6730 24828 6736 24880
rect 6788 24828 6794 24880
rect 7650 24828 7656 24880
rect 7708 24828 7714 24880
rect 8570 24828 8576 24880
rect 8628 24868 8634 24880
rect 9125 24871 9183 24877
rect 9125 24868 9137 24871
rect 8628 24840 9137 24868
rect 8628 24828 8634 24840
rect 9125 24837 9137 24840
rect 9171 24837 9183 24871
rect 9125 24831 9183 24837
rect 10778 24828 10784 24880
rect 10836 24828 10842 24880
rect 12710 24868 12716 24880
rect 11992 24840 12716 24868
rect 6822 24760 6828 24812
rect 6880 24760 6886 24812
rect 7024 24772 7972 24800
rect 7024 24741 7052 24772
rect 7944 24741 7972 24772
rect 8202 24760 8208 24812
rect 8260 24760 8266 24812
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8846 24800 8852 24812
rect 8352 24772 8852 24800
rect 8352 24760 8358 24772
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 10594 24800 10600 24812
rect 10258 24772 10600 24800
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10796 24800 10824 24828
rect 11992 24812 12020 24840
rect 12710 24828 12716 24840
rect 12768 24828 12774 24880
rect 13998 24828 14004 24880
rect 14056 24828 14062 24880
rect 16592 24868 16620 24896
rect 15672 24840 16620 24868
rect 16669 24871 16727 24877
rect 10796 24772 11560 24800
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24701 7067 24735
rect 7009 24695 7067 24701
rect 7745 24735 7803 24741
rect 7745 24701 7757 24735
rect 7791 24701 7803 24735
rect 7745 24695 7803 24701
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8110 24732 8116 24744
rect 7975 24704 8116 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 7760 24664 7788 24695
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 10870 24692 10876 24744
rect 10928 24692 10934 24744
rect 11532 24741 11560 24772
rect 11974 24760 11980 24812
rect 12032 24760 12038 24812
rect 12434 24760 12440 24812
rect 12492 24760 12498 24812
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24769 15439 24803
rect 15381 24763 15439 24769
rect 11517 24735 11575 24741
rect 11517 24701 11529 24735
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24701 13323 24735
rect 13265 24695 13323 24701
rect 8757 24667 8815 24673
rect 8757 24664 8769 24667
rect 7760 24636 8769 24664
rect 8757 24633 8769 24636
rect 8803 24633 8815 24667
rect 8757 24627 8815 24633
rect 11532 24608 11560 24695
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 12158 24664 12164 24676
rect 11931 24636 12164 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12158 24624 12164 24636
rect 12216 24624 12222 24676
rect 12802 24624 12808 24676
rect 12860 24664 12866 24676
rect 12989 24667 13047 24673
rect 12989 24664 13001 24667
rect 12860 24636 13001 24664
rect 12860 24624 12866 24636
rect 12989 24633 13001 24636
rect 13035 24633 13047 24667
rect 12989 24627 13047 24633
rect 7282 24556 7288 24608
rect 7340 24556 7346 24608
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 11330 24596 11336 24608
rect 9732 24568 11336 24596
rect 9732 24556 9738 24568
rect 11330 24556 11336 24568
rect 11388 24556 11394 24608
rect 11514 24556 11520 24608
rect 11572 24556 11578 24608
rect 12250 24556 12256 24608
rect 12308 24556 12314 24608
rect 13280 24596 13308 24695
rect 13538 24692 13544 24744
rect 13596 24692 13602 24744
rect 15396 24732 15424 24763
rect 15470 24760 15476 24812
rect 15528 24760 15534 24812
rect 15562 24760 15568 24812
rect 15620 24760 15626 24812
rect 15672 24732 15700 24840
rect 16669 24837 16681 24871
rect 16715 24868 16727 24871
rect 16850 24868 16856 24880
rect 16715 24840 16856 24868
rect 16715 24837 16727 24840
rect 16669 24831 16727 24837
rect 16850 24828 16856 24840
rect 16908 24868 16914 24880
rect 17586 24868 17592 24880
rect 16908 24840 17592 24868
rect 16908 24828 16914 24840
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 17770 24828 17776 24880
rect 17828 24828 17834 24880
rect 19444 24868 19472 24896
rect 19352 24840 19472 24868
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16758 24800 16764 24812
rect 16071 24772 16764 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 15396 24704 15700 24732
rect 15013 24667 15071 24673
rect 15013 24633 15025 24667
rect 15059 24664 15071 24667
rect 15102 24664 15108 24676
rect 15059 24636 15108 24664
rect 15059 24633 15071 24636
rect 15013 24627 15071 24633
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 13722 24596 13728 24608
rect 13280 24568 13728 24596
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 15764 24596 15792 24763
rect 16758 24760 16764 24772
rect 16816 24800 16822 24812
rect 17788 24800 17816 24828
rect 16816 24772 17816 24800
rect 16816 24760 16822 24772
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 19352 24800 19380 24840
rect 21174 24828 21180 24880
rect 21232 24868 21238 24880
rect 21232 24840 21680 24868
rect 21232 24828 21238 24840
rect 18196 24772 19380 24800
rect 18196 24760 18202 24772
rect 16117 24735 16175 24741
rect 16117 24701 16129 24735
rect 16163 24732 16175 24735
rect 16206 24732 16212 24744
rect 16163 24704 16212 24732
rect 16163 24701 16175 24704
rect 16117 24695 16175 24701
rect 16206 24692 16212 24704
rect 16264 24692 16270 24744
rect 17221 24735 17279 24741
rect 17221 24701 17233 24735
rect 17267 24701 17279 24735
rect 17221 24695 17279 24701
rect 16666 24624 16672 24676
rect 16724 24664 16730 24676
rect 16945 24667 17003 24673
rect 16945 24664 16957 24667
rect 16724 24636 16957 24664
rect 16724 24624 16730 24636
rect 16945 24633 16957 24636
rect 16991 24633 17003 24667
rect 17236 24664 17264 24695
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17681 24735 17739 24741
rect 17681 24732 17693 24735
rect 17368 24704 17693 24732
rect 17368 24692 17374 24704
rect 17681 24701 17693 24704
rect 17727 24701 17739 24735
rect 17681 24695 17739 24701
rect 17773 24735 17831 24741
rect 17773 24701 17785 24735
rect 17819 24732 17831 24735
rect 17819 24704 18276 24732
rect 17819 24701 17831 24704
rect 17773 24695 17831 24701
rect 17589 24667 17647 24673
rect 17236 24636 17356 24664
rect 16945 24627 17003 24633
rect 14700 24568 15792 24596
rect 14700 24556 14706 24568
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 17328 24596 17356 24636
rect 17589 24633 17601 24667
rect 17635 24664 17647 24667
rect 17788 24664 17816 24695
rect 17635 24636 17816 24664
rect 17635 24633 17647 24636
rect 17589 24627 17647 24633
rect 18138 24624 18144 24676
rect 18196 24624 18202 24676
rect 18248 24664 18276 24704
rect 19334 24692 19340 24744
rect 19392 24692 19398 24744
rect 19610 24692 19616 24744
rect 19668 24692 19674 24744
rect 20732 24664 20760 24786
rect 21358 24760 21364 24812
rect 21416 24760 21422 24812
rect 21652 24809 21680 24840
rect 21637 24803 21695 24809
rect 21637 24769 21649 24803
rect 21683 24769 21695 24803
rect 21637 24763 21695 24769
rect 21082 24692 21088 24744
rect 21140 24692 21146 24744
rect 21177 24667 21235 24673
rect 21177 24664 21189 24667
rect 18248 24636 19334 24664
rect 20732 24636 21189 24664
rect 18156 24596 18184 24624
rect 15896 24568 18184 24596
rect 15896 24556 15902 24568
rect 18230 24556 18236 24608
rect 18288 24556 18294 24608
rect 19306 24596 19334 24636
rect 21177 24633 21189 24636
rect 21223 24633 21235 24667
rect 21177 24627 21235 24633
rect 19794 24596 19800 24608
rect 19306 24568 19800 24596
rect 19794 24556 19800 24568
rect 19852 24556 19858 24608
rect 1104 24506 25852 24528
rect 1104 24454 4043 24506
rect 4095 24454 4107 24506
rect 4159 24454 4171 24506
rect 4223 24454 4235 24506
rect 4287 24454 4299 24506
rect 4351 24454 10230 24506
rect 10282 24454 10294 24506
rect 10346 24454 10358 24506
rect 10410 24454 10422 24506
rect 10474 24454 10486 24506
rect 10538 24454 16417 24506
rect 16469 24454 16481 24506
rect 16533 24454 16545 24506
rect 16597 24454 16609 24506
rect 16661 24454 16673 24506
rect 16725 24454 22604 24506
rect 22656 24454 22668 24506
rect 22720 24454 22732 24506
rect 22784 24454 22796 24506
rect 22848 24454 22860 24506
rect 22912 24454 25852 24506
rect 1104 24432 25852 24454
rect 7282 24352 7288 24404
rect 7340 24352 7346 24404
rect 8113 24395 8171 24401
rect 8113 24361 8125 24395
rect 8159 24392 8171 24395
rect 8662 24392 8668 24404
rect 8159 24364 8668 24392
rect 8159 24361 8171 24364
rect 8113 24355 8171 24361
rect 8662 24352 8668 24364
rect 8720 24352 8726 24404
rect 10413 24395 10471 24401
rect 10413 24361 10425 24395
rect 10459 24392 10471 24395
rect 10594 24392 10600 24404
rect 10459 24364 10600 24392
rect 10459 24361 10471 24364
rect 10413 24355 10471 24361
rect 10594 24352 10600 24364
rect 10652 24352 10658 24404
rect 11422 24392 11428 24404
rect 11072 24364 11428 24392
rect 7300 24188 7328 24352
rect 10229 24327 10287 24333
rect 10229 24293 10241 24327
rect 10275 24324 10287 24327
rect 11072 24324 11100 24364
rect 11422 24352 11428 24364
rect 11480 24392 11486 24404
rect 12158 24392 12164 24404
rect 11480 24364 12164 24392
rect 11480 24352 11486 24364
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 13538 24352 13544 24404
rect 13596 24392 13602 24404
rect 14093 24395 14151 24401
rect 14093 24392 14105 24395
rect 13596 24364 14105 24392
rect 13596 24352 13602 24364
rect 14093 24361 14105 24364
rect 14139 24361 14151 24395
rect 15289 24395 15347 24401
rect 14093 24355 14151 24361
rect 14200 24364 15148 24392
rect 13081 24327 13139 24333
rect 10275 24296 11100 24324
rect 11164 24296 11468 24324
rect 10275 24293 10287 24296
rect 10229 24287 10287 24293
rect 10321 24259 10379 24265
rect 10321 24225 10333 24259
rect 10367 24256 10379 24259
rect 10367 24228 10640 24256
rect 10367 24225 10379 24228
rect 10321 24219 10379 24225
rect 8297 24191 8355 24197
rect 8297 24188 8309 24191
rect 7300 24160 8309 24188
rect 8297 24157 8309 24160
rect 8343 24157 8355 24191
rect 8297 24151 8355 24157
rect 8386 24148 8392 24200
rect 8444 24188 8450 24200
rect 9122 24188 9128 24200
rect 8444 24160 9128 24188
rect 8444 24148 8450 24160
rect 9122 24148 9128 24160
rect 9180 24188 9186 24200
rect 10612 24197 10640 24228
rect 10597 24191 10655 24197
rect 9180 24160 10548 24188
rect 9180 24148 9186 24160
rect 934 24080 940 24132
rect 992 24120 998 24132
rect 1489 24123 1547 24129
rect 1489 24120 1501 24123
rect 992 24092 1501 24120
rect 992 24080 998 24092
rect 1489 24089 1501 24092
rect 1535 24089 1547 24123
rect 1489 24083 1547 24089
rect 9766 24080 9772 24132
rect 9824 24120 9830 24132
rect 9861 24123 9919 24129
rect 9861 24120 9873 24123
rect 9824 24092 9873 24120
rect 9824 24080 9830 24092
rect 9861 24089 9873 24092
rect 9907 24089 9919 24123
rect 10520 24120 10548 24160
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 11164 24120 11192 24296
rect 11238 24216 11244 24268
rect 11296 24256 11302 24268
rect 11333 24259 11391 24265
rect 11333 24256 11345 24259
rect 11296 24228 11345 24256
rect 11296 24216 11302 24228
rect 11333 24225 11345 24228
rect 11379 24225 11391 24259
rect 11440 24256 11468 24296
rect 13081 24293 13093 24327
rect 13127 24324 13139 24327
rect 14200 24324 14228 24364
rect 15120 24324 15148 24364
rect 15289 24361 15301 24395
rect 15335 24392 15347 24395
rect 15562 24392 15568 24404
rect 15335 24364 15568 24392
rect 15335 24361 15347 24364
rect 15289 24355 15347 24361
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 15838 24352 15844 24404
rect 15896 24352 15902 24404
rect 15930 24352 15936 24404
rect 15988 24352 15994 24404
rect 16850 24352 16856 24404
rect 16908 24392 16914 24404
rect 17497 24395 17555 24401
rect 17497 24392 17509 24395
rect 16908 24364 17509 24392
rect 16908 24352 16914 24364
rect 17497 24361 17509 24364
rect 17543 24361 17555 24395
rect 17497 24355 17555 24361
rect 20165 24395 20223 24401
rect 20165 24361 20177 24395
rect 20211 24392 20223 24395
rect 21358 24392 21364 24404
rect 20211 24364 21364 24392
rect 20211 24361 20223 24364
rect 20165 24355 20223 24361
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 15856 24324 15884 24352
rect 13127 24296 14228 24324
rect 14476 24296 15056 24324
rect 15120 24296 15884 24324
rect 15948 24324 15976 24352
rect 16485 24327 16543 24333
rect 15948 24296 16436 24324
rect 13127 24293 13139 24296
rect 13081 24287 13139 24293
rect 13372 24265 13400 24296
rect 13357 24259 13415 24265
rect 11440 24228 13308 24256
rect 11333 24219 11391 24225
rect 13280 24188 13308 24228
rect 13357 24225 13369 24259
rect 13403 24225 13415 24259
rect 14476 24256 14504 24296
rect 14921 24259 14979 24265
rect 14921 24256 14933 24259
rect 13357 24219 13415 24225
rect 13832 24228 14504 24256
rect 14568 24228 14933 24256
rect 13832 24188 13860 24228
rect 14568 24197 14596 24228
rect 14921 24225 14933 24228
rect 14967 24225 14979 24259
rect 14921 24219 14979 24225
rect 15028 24256 15056 24296
rect 15218 24256 15516 24264
rect 15028 24236 15516 24256
rect 15028 24228 15246 24236
rect 13280 24160 13860 24188
rect 13909 24191 13967 24197
rect 13909 24157 13921 24191
rect 13955 24188 13967 24191
rect 14369 24191 14427 24197
rect 14369 24188 14381 24191
rect 13955 24160 14381 24188
rect 13955 24157 13967 24160
rect 13909 24151 13967 24157
rect 14369 24157 14381 24160
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 10520 24092 11192 24120
rect 9861 24083 9919 24089
rect 1578 24012 1584 24064
rect 1636 24012 1642 24064
rect 9876 24052 9904 24083
rect 11330 24080 11336 24132
rect 11388 24120 11394 24132
rect 11609 24123 11667 24129
rect 11609 24120 11621 24123
rect 11388 24092 11621 24120
rect 11388 24080 11394 24092
rect 11609 24089 11621 24092
rect 11655 24089 11667 24123
rect 11609 24083 11667 24089
rect 12250 24080 12256 24132
rect 12308 24080 12314 24132
rect 14476 24064 14504 24151
rect 14642 24148 14648 24200
rect 14700 24188 14706 24200
rect 15028 24197 15056 24228
rect 14737 24191 14795 24197
rect 14737 24188 14749 24191
rect 14700 24160 14749 24188
rect 14700 24148 14706 24160
rect 14737 24157 14749 24160
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24157 15071 24191
rect 15013 24151 15071 24157
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24185 15255 24191
rect 15286 24185 15292 24200
rect 15243 24157 15292 24185
rect 15197 24151 15255 24157
rect 14844 24120 14872 24151
rect 15286 24148 15292 24157
rect 15344 24148 15350 24200
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15488 24188 15516 24236
rect 16408 24256 16436 24296
rect 16485 24293 16497 24327
rect 16531 24324 16543 24327
rect 17126 24324 17132 24336
rect 16531 24296 17132 24324
rect 16531 24293 16543 24296
rect 16485 24287 16543 24293
rect 17126 24284 17132 24296
rect 17184 24284 17190 24336
rect 20070 24284 20076 24336
rect 20128 24324 20134 24336
rect 20625 24327 20683 24333
rect 20625 24324 20637 24327
rect 20128 24296 20637 24324
rect 20128 24284 20134 24296
rect 20625 24293 20637 24296
rect 20671 24293 20683 24327
rect 20625 24287 20683 24293
rect 16577 24259 16635 24265
rect 16577 24256 16589 24259
rect 16408 24228 16589 24256
rect 16577 24225 16589 24228
rect 16623 24225 16635 24259
rect 16942 24256 16948 24268
rect 16577 24219 16635 24225
rect 16684 24228 16948 24256
rect 15427 24160 15516 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15654 24148 15660 24200
rect 15712 24148 15718 24200
rect 16114 24148 16120 24200
rect 16172 24188 16178 24200
rect 16684 24197 16712 24228
rect 16942 24216 16948 24228
rect 17000 24256 17006 24268
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 17000 24228 17601 24256
rect 17000 24216 17006 24228
rect 17589 24225 17601 24228
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 20809 24259 20867 24265
rect 20809 24225 20821 24259
rect 20855 24256 20867 24259
rect 20855 24228 21680 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 16172 24160 16405 24188
rect 16172 24148 16178 24160
rect 16393 24157 16405 24160
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 17126 24188 17132 24200
rect 16899 24160 17132 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 16408 24120 16436 24151
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17037 24123 17095 24129
rect 17037 24120 17049 24123
rect 14844 24092 16160 24120
rect 16408 24092 17049 24120
rect 11514 24052 11520 24064
rect 9876 24024 11520 24052
rect 11514 24012 11520 24024
rect 11572 24052 11578 24064
rect 14366 24052 14372 24064
rect 11572 24024 14372 24052
rect 11572 24012 11578 24024
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 15470 24052 15476 24064
rect 14516 24024 15476 24052
rect 14516 24012 14522 24024
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 16132 24061 16160 24092
rect 17037 24089 17049 24092
rect 17083 24120 17095 24123
rect 17328 24120 17356 24151
rect 17402 24148 17408 24200
rect 17460 24148 17466 24200
rect 17494 24148 17500 24200
rect 17552 24188 17558 24200
rect 19518 24188 19524 24200
rect 17552 24160 19524 24188
rect 17552 24148 17558 24160
rect 19518 24148 19524 24160
rect 19576 24188 19582 24200
rect 19705 24191 19763 24197
rect 19705 24188 19717 24191
rect 19576 24160 19717 24188
rect 19576 24148 19582 24160
rect 19705 24157 19717 24160
rect 19751 24188 19763 24191
rect 19978 24188 19984 24200
rect 19751 24160 19984 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 19978 24148 19984 24160
rect 20036 24188 20042 24200
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 20036 24160 20361 24188
rect 20036 24148 20042 24160
rect 20349 24157 20361 24160
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 21358 24148 21364 24200
rect 21416 24148 21422 24200
rect 21652 24197 21680 24228
rect 21637 24191 21695 24197
rect 21637 24157 21649 24191
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 18230 24120 18236 24132
rect 17083 24092 18236 24120
rect 17083 24089 17095 24092
rect 17037 24083 17095 24089
rect 18230 24080 18236 24092
rect 18288 24080 18294 24132
rect 22002 24120 22008 24132
rect 21192 24092 22008 24120
rect 16117 24055 16175 24061
rect 16117 24021 16129 24055
rect 16163 24021 16175 24055
rect 16117 24015 16175 24021
rect 16206 24012 16212 24064
rect 16264 24012 16270 24064
rect 16942 24012 16948 24064
rect 17000 24052 17006 24064
rect 21192 24061 21220 24092
rect 22002 24080 22008 24092
rect 22060 24080 22066 24132
rect 17221 24055 17279 24061
rect 17221 24052 17233 24055
rect 17000 24024 17233 24052
rect 17000 24012 17006 24024
rect 17221 24021 17233 24024
rect 17267 24021 17279 24055
rect 17221 24015 17279 24021
rect 21177 24055 21235 24061
rect 21177 24021 21189 24055
rect 21223 24021 21235 24055
rect 21177 24015 21235 24021
rect 21450 24012 21456 24064
rect 21508 24012 21514 24064
rect 25406 24012 25412 24064
rect 25464 24012 25470 24064
rect 1104 23962 25852 23984
rect 1104 23910 4703 23962
rect 4755 23910 4767 23962
rect 4819 23910 4831 23962
rect 4883 23910 4895 23962
rect 4947 23910 4959 23962
rect 5011 23910 10890 23962
rect 10942 23910 10954 23962
rect 11006 23910 11018 23962
rect 11070 23910 11082 23962
rect 11134 23910 11146 23962
rect 11198 23910 17077 23962
rect 17129 23910 17141 23962
rect 17193 23910 17205 23962
rect 17257 23910 17269 23962
rect 17321 23910 17333 23962
rect 17385 23910 23264 23962
rect 23316 23910 23328 23962
rect 23380 23910 23392 23962
rect 23444 23910 23456 23962
rect 23508 23910 23520 23962
rect 23572 23910 25852 23962
rect 1104 23888 25852 23910
rect 1578 23808 1584 23860
rect 1636 23808 1642 23860
rect 9401 23851 9459 23857
rect 9401 23817 9413 23851
rect 9447 23848 9459 23851
rect 9628 23848 9634 23860
rect 9447 23820 9634 23848
rect 9447 23817 9459 23820
rect 9401 23811 9459 23817
rect 9628 23808 9634 23820
rect 9686 23808 9692 23860
rect 9766 23808 9772 23860
rect 9824 23808 9830 23860
rect 12253 23851 12311 23857
rect 12253 23817 12265 23851
rect 12299 23848 12311 23851
rect 12434 23848 12440 23860
rect 12299 23820 12440 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 12434 23808 12440 23820
rect 12492 23808 12498 23860
rect 13725 23851 13783 23857
rect 13725 23817 13737 23851
rect 13771 23848 13783 23851
rect 13998 23848 14004 23860
rect 13771 23820 14004 23848
rect 13771 23817 13783 23820
rect 13725 23811 13783 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15841 23851 15899 23857
rect 15841 23848 15853 23851
rect 15712 23820 15853 23848
rect 15712 23808 15718 23820
rect 15841 23817 15853 23820
rect 15887 23817 15899 23851
rect 15841 23811 15899 23817
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 16117 23851 16175 23857
rect 16117 23848 16129 23851
rect 15988 23820 16129 23848
rect 15988 23808 15994 23820
rect 16117 23817 16129 23820
rect 16163 23817 16175 23851
rect 16117 23811 16175 23817
rect 16298 23808 16304 23860
rect 16356 23848 16362 23860
rect 17037 23851 17095 23857
rect 17037 23848 17049 23851
rect 16356 23820 17049 23848
rect 16356 23808 16362 23820
rect 17037 23817 17049 23820
rect 17083 23817 17095 23851
rect 17037 23811 17095 23817
rect 19610 23808 19616 23860
rect 19668 23848 19674 23860
rect 20165 23851 20223 23857
rect 20165 23848 20177 23851
rect 19668 23820 20177 23848
rect 19668 23808 19674 23820
rect 20165 23817 20177 23820
rect 20211 23817 20223 23851
rect 20165 23811 20223 23817
rect 20901 23851 20959 23857
rect 20901 23817 20913 23851
rect 20947 23848 20959 23851
rect 21358 23848 21364 23860
rect 20947 23820 21364 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 21450 23808 21456 23860
rect 21508 23848 21514 23860
rect 21508 23820 22416 23848
rect 21508 23808 21514 23820
rect 1394 23672 1400 23724
rect 1452 23672 1458 23724
rect 1596 23644 1624 23808
rect 9784 23780 9812 23808
rect 2746 23752 9812 23780
rect 2746 23644 2774 23752
rect 11790 23740 11796 23792
rect 11848 23780 11854 23792
rect 11974 23780 11980 23792
rect 11848 23752 11980 23780
rect 11848 23740 11854 23752
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 13814 23740 13820 23792
rect 13872 23740 13878 23792
rect 16758 23780 16764 23792
rect 14016 23752 16436 23780
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 5316 23684 5549 23712
rect 5316 23672 5322 23684
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 5537 23675 5595 23681
rect 6178 23672 6184 23724
rect 6236 23712 6242 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 6236 23684 6561 23712
rect 6236 23672 6242 23684
rect 6549 23681 6561 23684
rect 6595 23681 6607 23715
rect 8205 23715 8263 23721
rect 8205 23712 8217 23715
rect 6549 23675 6607 23681
rect 6932 23684 8217 23712
rect 1596 23616 2774 23644
rect 5718 23604 5724 23656
rect 5776 23644 5782 23656
rect 5813 23647 5871 23653
rect 5813 23644 5825 23647
rect 5776 23616 5825 23644
rect 5776 23604 5782 23616
rect 5813 23613 5825 23616
rect 5859 23613 5871 23647
rect 5813 23607 5871 23613
rect 5994 23604 6000 23656
rect 6052 23644 6058 23656
rect 6457 23647 6515 23653
rect 6457 23644 6469 23647
rect 6052 23616 6469 23644
rect 6052 23604 6058 23616
rect 6457 23613 6469 23616
rect 6503 23613 6515 23647
rect 6457 23607 6515 23613
rect 1578 23536 1584 23588
rect 1636 23536 1642 23588
rect 5353 23579 5411 23585
rect 5353 23545 5365 23579
rect 5399 23576 5411 23579
rect 5902 23576 5908 23588
rect 5399 23548 5908 23576
rect 5399 23545 5411 23548
rect 5353 23539 5411 23545
rect 5902 23536 5908 23548
rect 5960 23536 5966 23588
rect 6932 23585 6960 23684
rect 8205 23681 8217 23684
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 8386 23672 8392 23724
rect 8444 23672 8450 23724
rect 9490 23672 9496 23724
rect 9548 23718 9554 23724
rect 9631 23718 9689 23721
rect 9548 23715 9689 23718
rect 9548 23690 9643 23715
rect 9548 23672 9554 23690
rect 9631 23681 9643 23690
rect 9677 23681 9689 23715
rect 9631 23675 9689 23681
rect 9766 23672 9772 23724
rect 9824 23672 9830 23724
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23687 10272 23715
rect 10091 23681 10103 23687
rect 10045 23675 10103 23681
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23644 8355 23647
rect 9876 23644 9904 23675
rect 8343 23616 9904 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 10134 23604 10140 23656
rect 10192 23644 10198 23656
rect 10244 23644 10272 23687
rect 10318 23672 10324 23724
rect 10376 23672 10382 23724
rect 13832 23712 13860 23740
rect 13909 23715 13967 23721
rect 13909 23712 13921 23715
rect 13832 23684 13921 23712
rect 13909 23681 13921 23684
rect 13955 23681 13967 23715
rect 13909 23675 13967 23681
rect 10192 23616 10272 23644
rect 10192 23604 10198 23616
rect 10502 23604 10508 23656
rect 10560 23644 10566 23656
rect 14016 23644 14044 23752
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 15749 23715 15807 23721
rect 15749 23712 15761 23715
rect 15712 23684 15761 23712
rect 15712 23672 15718 23684
rect 15749 23681 15761 23684
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 10560 23616 14044 23644
rect 15956 23644 15984 23675
rect 16022 23672 16028 23724
rect 16080 23721 16086 23724
rect 16080 23712 16089 23721
rect 16209 23715 16267 23721
rect 16080 23684 16125 23712
rect 16080 23675 16089 23684
rect 16209 23681 16221 23715
rect 16255 23712 16267 23715
rect 16255 23684 16344 23712
rect 16255 23681 16267 23684
rect 16209 23675 16267 23681
rect 16080 23672 16086 23675
rect 15956 23616 16068 23644
rect 10560 23604 10566 23616
rect 16040 23588 16068 23616
rect 6917 23579 6975 23585
rect 6917 23545 6929 23579
rect 6963 23545 6975 23579
rect 6917 23539 6975 23545
rect 10042 23536 10048 23588
rect 10100 23576 10106 23588
rect 10410 23576 10416 23588
rect 10100 23548 10416 23576
rect 10100 23536 10106 23548
rect 10410 23536 10416 23548
rect 10468 23536 10474 23588
rect 12161 23579 12219 23585
rect 12161 23545 12173 23579
rect 12207 23576 12219 23579
rect 12250 23576 12256 23588
rect 12207 23548 12256 23576
rect 12207 23545 12219 23548
rect 12161 23539 12219 23545
rect 12250 23536 12256 23548
rect 12308 23576 12314 23588
rect 12802 23576 12808 23588
rect 12308 23548 12808 23576
rect 12308 23536 12314 23548
rect 12802 23536 12808 23548
rect 12860 23536 12866 23588
rect 16022 23536 16028 23588
rect 16080 23576 16086 23588
rect 16316 23576 16344 23684
rect 16408 23644 16436 23752
rect 16684 23752 16764 23780
rect 16684 23721 16712 23752
rect 16758 23740 16764 23752
rect 16816 23740 16822 23792
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 19392 23752 21864 23780
rect 19392 23740 19398 23752
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23712 16911 23715
rect 17586 23712 17592 23724
rect 16899 23684 17592 23712
rect 16899 23681 16911 23684
rect 16853 23675 16911 23681
rect 17586 23672 17592 23684
rect 17644 23672 17650 23724
rect 19794 23712 19800 23724
rect 19306 23684 19800 23712
rect 19306 23644 19334 23684
rect 19794 23672 19800 23684
rect 19852 23672 19858 23724
rect 19978 23672 19984 23724
rect 20036 23672 20042 23724
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23681 20407 23715
rect 20349 23675 20407 23681
rect 16408 23616 19334 23644
rect 20364 23644 20392 23675
rect 20714 23672 20720 23724
rect 20772 23672 20778 23724
rect 21266 23672 21272 23724
rect 21324 23672 21330 23724
rect 21836 23721 21864 23752
rect 22002 23740 22008 23792
rect 22060 23780 22066 23792
rect 22097 23783 22155 23789
rect 22097 23780 22109 23783
rect 22060 23752 22109 23780
rect 22060 23740 22066 23752
rect 22097 23749 22109 23752
rect 22143 23749 22155 23783
rect 22388 23780 22416 23820
rect 22388 23752 22586 23780
rect 22097 23743 22155 23749
rect 21821 23715 21879 23721
rect 21821 23681 21833 23715
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 25317 23715 25375 23721
rect 25317 23681 25329 23715
rect 25363 23712 25375 23715
rect 25363 23684 25820 23712
rect 25363 23681 25375 23684
rect 25317 23675 25375 23681
rect 20898 23644 20904 23656
rect 20364 23616 20904 23644
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23613 21419 23647
rect 21361 23607 21419 23613
rect 16080 23548 16344 23576
rect 16080 23536 16086 23548
rect 16390 23536 16396 23588
rect 16448 23576 16454 23588
rect 19518 23576 19524 23588
rect 16448 23548 19524 23576
rect 16448 23536 16454 23548
rect 19518 23536 19524 23548
rect 19576 23536 19582 23588
rect 21376 23576 21404 23607
rect 21542 23604 21548 23656
rect 21600 23604 21606 23656
rect 22186 23644 22192 23656
rect 21744 23616 22192 23644
rect 21744 23576 21772 23616
rect 22186 23604 22192 23616
rect 22244 23644 22250 23656
rect 25590 23644 25596 23656
rect 22244 23616 25596 23644
rect 22244 23604 22250 23616
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 21376 23548 21772 23576
rect 25792 23520 25820 23684
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 5721 23511 5779 23517
rect 5721 23508 5733 23511
rect 5592 23480 5733 23508
rect 5592 23468 5598 23480
rect 5721 23477 5733 23480
rect 5767 23508 5779 23511
rect 6822 23508 6828 23520
rect 5767 23480 6828 23508
rect 5767 23477 5779 23480
rect 5721 23471 5779 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 8662 23468 8668 23520
rect 8720 23508 8726 23520
rect 9766 23508 9772 23520
rect 8720 23480 9772 23508
rect 8720 23468 8726 23480
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 9950 23468 9956 23520
rect 10008 23508 10014 23520
rect 10137 23511 10195 23517
rect 10137 23508 10149 23511
rect 10008 23480 10149 23508
rect 10008 23468 10014 23480
rect 10137 23477 10149 23480
rect 10183 23477 10195 23511
rect 10137 23471 10195 23477
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 16942 23508 16948 23520
rect 16899 23480 16948 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 20533 23511 20591 23517
rect 20533 23477 20545 23511
rect 20579 23508 20591 23511
rect 20990 23508 20996 23520
rect 20579 23480 20996 23508
rect 20579 23477 20591 23480
rect 20533 23471 20591 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21542 23468 21548 23520
rect 21600 23508 21606 23520
rect 21818 23508 21824 23520
rect 21600 23480 21824 23508
rect 21600 23468 21606 23480
rect 21818 23468 21824 23480
rect 21876 23468 21882 23520
rect 23569 23511 23627 23517
rect 23569 23477 23581 23511
rect 23615 23508 23627 23511
rect 23750 23508 23756 23520
rect 23615 23480 23756 23508
rect 23615 23477 23627 23480
rect 23569 23471 23627 23477
rect 23750 23468 23756 23480
rect 23808 23508 23814 23520
rect 24302 23508 24308 23520
rect 23808 23480 24308 23508
rect 23808 23468 23814 23480
rect 24302 23468 24308 23480
rect 24360 23468 24366 23520
rect 25498 23468 25504 23520
rect 25556 23468 25562 23520
rect 25774 23468 25780 23520
rect 25832 23468 25838 23520
rect 1104 23418 25852 23440
rect 1104 23366 4043 23418
rect 4095 23366 4107 23418
rect 4159 23366 4171 23418
rect 4223 23366 4235 23418
rect 4287 23366 4299 23418
rect 4351 23366 10230 23418
rect 10282 23366 10294 23418
rect 10346 23366 10358 23418
rect 10410 23366 10422 23418
rect 10474 23366 10486 23418
rect 10538 23366 16417 23418
rect 16469 23366 16481 23418
rect 16533 23366 16545 23418
rect 16597 23366 16609 23418
rect 16661 23366 16673 23418
rect 16725 23366 22604 23418
rect 22656 23366 22668 23418
rect 22720 23366 22732 23418
rect 22784 23366 22796 23418
rect 22848 23366 22860 23418
rect 22912 23366 25852 23418
rect 1104 23344 25852 23366
rect 6822 23264 6828 23316
rect 6880 23304 6886 23316
rect 6880 23276 9076 23304
rect 6880 23264 6886 23276
rect 3602 23196 3608 23248
rect 3660 23236 3666 23248
rect 4525 23239 4583 23245
rect 4525 23236 4537 23239
rect 3660 23208 4537 23236
rect 3660 23196 3666 23208
rect 4525 23205 4537 23208
rect 4571 23205 4583 23239
rect 4525 23199 4583 23205
rect 5169 23239 5227 23245
rect 5169 23205 5181 23239
rect 5215 23236 5227 23239
rect 5215 23208 5396 23236
rect 5215 23205 5227 23208
rect 5169 23199 5227 23205
rect 4540 23168 4568 23199
rect 4801 23171 4859 23177
rect 4801 23168 4813 23171
rect 4540 23140 4813 23168
rect 4801 23137 4813 23140
rect 4847 23137 4859 23171
rect 4801 23131 4859 23137
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 5368 23100 5396 23208
rect 6012 23208 7604 23236
rect 5534 23100 5540 23112
rect 4295 23072 5396 23100
rect 5498 23072 5540 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 5368 23032 5396 23072
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5718 23100 5724 23112
rect 5675 23072 5724 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5810 23060 5816 23112
rect 5868 23060 5874 23112
rect 5902 23060 5908 23112
rect 5960 23060 5966 23112
rect 6012 23032 6040 23208
rect 7576 23180 7604 23208
rect 6362 23128 6368 23180
rect 6420 23128 6426 23180
rect 6638 23128 6644 23180
rect 6696 23128 6702 23180
rect 7558 23128 7564 23180
rect 7616 23128 7622 23180
rect 8846 23128 8852 23180
rect 8904 23168 8910 23180
rect 8941 23171 8999 23177
rect 8941 23168 8953 23171
rect 8904 23140 8953 23168
rect 8904 23128 8910 23140
rect 8941 23137 8953 23140
rect 8987 23137 8999 23171
rect 9048 23168 9076 23276
rect 9766 23264 9772 23316
rect 9824 23304 9830 23316
rect 14458 23304 14464 23316
rect 9824 23276 14464 23304
rect 9824 23264 9830 23276
rect 14458 23264 14464 23276
rect 14516 23264 14522 23316
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 15930 23304 15936 23316
rect 15712 23276 15936 23304
rect 15712 23264 15718 23276
rect 15930 23264 15936 23276
rect 15988 23304 15994 23316
rect 16942 23304 16948 23316
rect 15988 23276 16948 23304
rect 15988 23264 15994 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 20349 23307 20407 23313
rect 20349 23273 20361 23307
rect 20395 23304 20407 23307
rect 20714 23304 20720 23316
rect 20395 23276 20720 23304
rect 20395 23273 20407 23276
rect 20349 23267 20407 23273
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 20898 23264 20904 23316
rect 20956 23264 20962 23316
rect 16206 23196 16212 23248
rect 16264 23236 16270 23248
rect 16264 23208 16988 23236
rect 16264 23196 16270 23208
rect 9582 23168 9588 23180
rect 9048 23140 9588 23168
rect 8941 23131 8999 23137
rect 9582 23128 9588 23140
rect 9640 23168 9646 23180
rect 10965 23171 11023 23177
rect 10965 23168 10977 23171
rect 9640 23140 10977 23168
rect 9640 23128 9646 23140
rect 10965 23137 10977 23140
rect 11011 23137 11023 23171
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 10965 23131 11023 23137
rect 12360 23140 12817 23168
rect 6086 23060 6092 23112
rect 6144 23100 6150 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 6144 23072 6285 23100
rect 6144 23060 6150 23072
rect 6273 23069 6285 23072
rect 6319 23100 6331 23103
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6319 23072 6745 23100
rect 6319 23069 6331 23072
rect 6273 23063 6331 23069
rect 6733 23069 6745 23072
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23100 7067 23103
rect 7650 23100 7656 23112
rect 7055 23072 7656 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 12360 23109 12388 23140
rect 12805 23137 12817 23140
rect 12851 23137 12863 23171
rect 12805 23131 12863 23137
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23069 12587 23103
rect 12529 23063 12587 23069
rect 5368 23004 6040 23032
rect 6178 22992 6184 23044
rect 6236 23032 6242 23044
rect 6917 23035 6975 23041
rect 6917 23032 6929 23035
rect 6236 23004 6929 23032
rect 6236 22992 6242 23004
rect 6917 23001 6929 23004
rect 6963 23001 6975 23035
rect 6917 22995 6975 23001
rect 9214 22992 9220 23044
rect 9272 22992 9278 23044
rect 9950 22992 9956 23044
rect 10008 22992 10014 23044
rect 11330 22992 11336 23044
rect 11388 23032 11394 23044
rect 12544 23032 12572 23063
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 14274 23060 14280 23112
rect 14332 23060 14338 23112
rect 14550 23060 14556 23112
rect 14608 23060 14614 23112
rect 16114 23060 16120 23112
rect 16172 23100 16178 23112
rect 16298 23100 16304 23112
rect 16172 23072 16304 23100
rect 16172 23060 16178 23072
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23100 16727 23103
rect 16758 23100 16764 23112
rect 16715 23072 16764 23100
rect 16715 23069 16727 23072
rect 16669 23063 16727 23069
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 16960 23109 16988 23208
rect 19518 23196 19524 23248
rect 19576 23236 19582 23248
rect 20070 23236 20076 23248
rect 19576 23208 20076 23236
rect 19576 23196 19582 23208
rect 20070 23196 20076 23208
rect 20128 23236 20134 23248
rect 20165 23239 20223 23245
rect 20165 23236 20177 23239
rect 20128 23208 20177 23236
rect 20128 23196 20134 23208
rect 20165 23205 20177 23208
rect 20211 23205 20223 23239
rect 20165 23199 20223 23205
rect 19245 23171 19303 23177
rect 19245 23137 19257 23171
rect 19291 23168 19303 23171
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 19291 23140 19901 23168
rect 19291 23137 19303 23140
rect 19245 23131 19303 23137
rect 19889 23137 19901 23140
rect 19935 23168 19947 23171
rect 19978 23168 19984 23180
rect 19935 23140 19984 23168
rect 19935 23137 19947 23140
rect 19889 23131 19947 23137
rect 19978 23128 19984 23140
rect 20036 23128 20042 23180
rect 16945 23103 17003 23109
rect 16945 23069 16957 23103
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 17037 23103 17095 23109
rect 17037 23069 17049 23103
rect 17083 23100 17095 23103
rect 17402 23100 17408 23112
rect 17083 23072 17408 23100
rect 17083 23069 17095 23072
rect 17037 23063 17095 23069
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23100 17555 23103
rect 17543 23072 17724 23100
rect 17543 23069 17555 23072
rect 17497 23063 17555 23069
rect 14568 23032 14596 23060
rect 11388 23004 14596 23032
rect 16776 23032 16804 23060
rect 17221 23035 17279 23041
rect 17221 23032 17233 23035
rect 16776 23004 17233 23032
rect 11388 22992 11394 23004
rect 17221 23001 17233 23004
rect 17267 23001 17279 23035
rect 17589 23035 17647 23041
rect 17589 23032 17601 23035
rect 17221 22995 17279 23001
rect 17328 23004 17601 23032
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 4709 22967 4767 22973
rect 4709 22964 4721 22967
rect 4672 22936 4721 22964
rect 4672 22924 4678 22936
rect 4709 22933 4721 22936
rect 4755 22933 4767 22967
rect 4709 22927 4767 22933
rect 5258 22924 5264 22976
rect 5316 22924 5322 22976
rect 5353 22967 5411 22973
rect 5353 22933 5365 22967
rect 5399 22964 5411 22967
rect 6822 22964 6828 22976
rect 5399 22936 6828 22964
rect 5399 22933 5411 22936
rect 5353 22927 5411 22933
rect 6822 22924 6828 22936
rect 6880 22924 6886 22976
rect 7098 22924 7104 22976
rect 7156 22924 7162 22976
rect 7282 22924 7288 22976
rect 7340 22924 7346 22976
rect 12158 22924 12164 22976
rect 12216 22924 12222 22976
rect 14090 22924 14096 22976
rect 14148 22924 14154 22976
rect 16298 22924 16304 22976
rect 16356 22964 16362 22976
rect 16485 22967 16543 22973
rect 16485 22964 16497 22967
rect 16356 22936 16497 22964
rect 16356 22924 16362 22936
rect 16485 22933 16497 22936
rect 16531 22933 16543 22967
rect 16485 22927 16543 22933
rect 16853 22967 16911 22973
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 17328 22964 17356 23004
rect 17589 23001 17601 23004
rect 17635 23001 17647 23035
rect 17589 22995 17647 23001
rect 16899 22936 17356 22964
rect 17405 22967 17463 22973
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 17405 22933 17417 22967
rect 17451 22964 17463 22967
rect 17494 22964 17500 22976
rect 17451 22936 17500 22964
rect 17451 22933 17463 22936
rect 17405 22927 17463 22933
rect 17494 22924 17500 22936
rect 17552 22964 17558 22976
rect 17696 22964 17724 23072
rect 17552 22936 17724 22964
rect 17552 22924 17558 22936
rect 19702 22924 19708 22976
rect 19760 22924 19766 22976
rect 20180 22964 20208 23199
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 21453 23171 21511 23177
rect 21453 23168 21465 23171
rect 20680 23140 21465 23168
rect 20680 23128 20686 23140
rect 21453 23137 21465 23140
rect 21499 23137 21511 23171
rect 21453 23131 21511 23137
rect 21821 23171 21879 23177
rect 21821 23137 21833 23171
rect 21867 23168 21879 23171
rect 21910 23168 21916 23180
rect 21867 23140 21916 23168
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 21910 23128 21916 23140
rect 21968 23128 21974 23180
rect 20530 23060 20536 23112
rect 20588 23060 20594 23112
rect 20717 22967 20775 22973
rect 20717 22964 20729 22967
rect 20180 22936 20729 22964
rect 20717 22933 20729 22936
rect 20763 22933 20775 22967
rect 20717 22927 20775 22933
rect 21266 22924 21272 22976
rect 21324 22924 21330 22976
rect 21361 22967 21419 22973
rect 21361 22933 21373 22967
rect 21407 22964 21419 22967
rect 22373 22967 22431 22973
rect 22373 22964 22385 22967
rect 21407 22936 22385 22964
rect 21407 22933 21419 22936
rect 21361 22927 21419 22933
rect 22373 22933 22385 22936
rect 22419 22933 22431 22967
rect 22373 22927 22431 22933
rect 1104 22874 25852 22896
rect 1104 22822 4703 22874
rect 4755 22822 4767 22874
rect 4819 22822 4831 22874
rect 4883 22822 4895 22874
rect 4947 22822 4959 22874
rect 5011 22822 10890 22874
rect 10942 22822 10954 22874
rect 11006 22822 11018 22874
rect 11070 22822 11082 22874
rect 11134 22822 11146 22874
rect 11198 22822 17077 22874
rect 17129 22822 17141 22874
rect 17193 22822 17205 22874
rect 17257 22822 17269 22874
rect 17321 22822 17333 22874
rect 17385 22822 23264 22874
rect 23316 22822 23328 22874
rect 23380 22822 23392 22874
rect 23444 22822 23456 22874
rect 23508 22822 23520 22874
rect 23572 22822 25852 22874
rect 1104 22800 25852 22822
rect 3050 22720 3056 22772
rect 3108 22760 3114 22772
rect 3329 22763 3387 22769
rect 3329 22760 3341 22763
rect 3108 22732 3341 22760
rect 3108 22720 3114 22732
rect 3329 22729 3341 22732
rect 3375 22760 3387 22763
rect 3694 22760 3700 22772
rect 3375 22732 3700 22760
rect 3375 22729 3387 22732
rect 3329 22723 3387 22729
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 6089 22763 6147 22769
rect 6089 22760 6101 22763
rect 5776 22732 6101 22760
rect 5776 22720 5782 22732
rect 6089 22729 6101 22732
rect 6135 22729 6147 22763
rect 6089 22723 6147 22729
rect 6638 22720 6644 22772
rect 6696 22760 6702 22772
rect 7561 22763 7619 22769
rect 7561 22760 7573 22763
rect 6696 22732 7573 22760
rect 6696 22720 6702 22732
rect 7561 22729 7573 22732
rect 7607 22729 7619 22763
rect 8202 22760 8208 22772
rect 7561 22723 7619 22729
rect 7668 22732 8208 22760
rect 3786 22652 3792 22704
rect 3844 22692 3850 22704
rect 3844 22664 4752 22692
rect 3844 22652 3850 22664
rect 1489 22627 1547 22633
rect 1489 22593 1501 22627
rect 1535 22624 1547 22627
rect 2498 22624 2504 22636
rect 1535 22596 2504 22624
rect 1535 22593 1547 22596
rect 1489 22587 1547 22593
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 4724 22633 4752 22664
rect 7006 22652 7012 22704
rect 7064 22692 7070 22704
rect 7668 22692 7696 22732
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 8389 22763 8447 22769
rect 8389 22729 8401 22763
rect 8435 22760 8447 22763
rect 9214 22760 9220 22772
rect 8435 22732 9220 22760
rect 8435 22729 8447 22732
rect 8389 22723 8447 22729
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 10229 22763 10287 22769
rect 10229 22760 10241 22763
rect 10192 22732 10241 22760
rect 10192 22720 10198 22732
rect 10229 22729 10241 22732
rect 10275 22729 10287 22763
rect 10229 22723 10287 22729
rect 11330 22720 11336 22772
rect 11388 22720 11394 22772
rect 12158 22760 12164 22772
rect 11900 22732 12164 22760
rect 11348 22692 11376 22720
rect 11900 22701 11928 22732
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 12618 22720 12624 22772
rect 12676 22760 12682 22772
rect 13725 22763 13783 22769
rect 13725 22760 13737 22763
rect 12676 22732 13737 22760
rect 12676 22720 12682 22732
rect 13725 22729 13737 22732
rect 13771 22729 13783 22763
rect 13725 22723 13783 22729
rect 14182 22720 14188 22772
rect 14240 22720 14246 22772
rect 14274 22720 14280 22772
rect 14332 22760 14338 22772
rect 15013 22763 15071 22769
rect 15013 22760 15025 22763
rect 14332 22732 15025 22760
rect 14332 22720 14338 22732
rect 15013 22729 15025 22732
rect 15059 22729 15071 22763
rect 17310 22760 17316 22772
rect 15013 22723 15071 22729
rect 16040 22732 17316 22760
rect 7064 22664 7696 22692
rect 7064 22652 7070 22664
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22624 2651 22627
rect 3421 22627 3479 22633
rect 2639 22596 2774 22624
rect 2639 22593 2651 22596
rect 2593 22587 2651 22593
rect 2746 22488 2774 22596
rect 3421 22593 3433 22627
rect 3467 22624 3479 22627
rect 4433 22627 4491 22633
rect 4433 22624 4445 22627
rect 3467 22596 4445 22624
rect 3467 22593 3479 22596
rect 3421 22587 3479 22593
rect 4433 22593 4445 22596
rect 4479 22593 4491 22627
rect 4433 22587 4491 22593
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22593 4767 22627
rect 4709 22587 4767 22593
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5997 22627 6055 22633
rect 5997 22624 6009 22627
rect 5132 22596 6009 22624
rect 5132 22584 5138 22596
rect 5997 22593 6009 22596
rect 6043 22593 6055 22627
rect 5997 22587 6055 22593
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 7190 22624 7196 22636
rect 6687 22596 7196 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 7515 22596 7604 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 7576 22568 7604 22596
rect 3513 22559 3571 22565
rect 3513 22525 3525 22559
rect 3559 22525 3571 22559
rect 3513 22519 3571 22525
rect 2961 22491 3019 22497
rect 2961 22488 2973 22491
rect 2746 22460 2973 22488
rect 2961 22457 2973 22460
rect 3007 22457 3019 22491
rect 3528 22488 3556 22519
rect 3602 22516 3608 22568
rect 3660 22556 3666 22568
rect 3789 22559 3847 22565
rect 3789 22556 3801 22559
rect 3660 22528 3801 22556
rect 3660 22516 3666 22528
rect 3789 22525 3801 22528
rect 3835 22525 3847 22559
rect 3789 22519 3847 22525
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22556 5411 22559
rect 5534 22556 5540 22568
rect 5399 22528 5540 22556
rect 5399 22525 5411 22528
rect 5353 22519 5411 22525
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 5718 22516 5724 22568
rect 5776 22556 5782 22568
rect 5813 22559 5871 22565
rect 5813 22556 5825 22559
rect 5776 22528 5825 22556
rect 5776 22516 5782 22528
rect 5813 22525 5825 22528
rect 5859 22556 5871 22559
rect 6178 22556 6184 22568
rect 5859 22528 6184 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 6178 22516 6184 22528
rect 6236 22516 6242 22568
rect 6733 22559 6791 22565
rect 6733 22525 6745 22559
rect 6779 22556 6791 22559
rect 6914 22556 6920 22568
rect 6779 22528 6920 22556
rect 6779 22525 6791 22528
rect 6733 22519 6791 22525
rect 6914 22516 6920 22528
rect 6972 22516 6978 22568
rect 7558 22516 7564 22568
rect 7616 22516 7622 22568
rect 7668 22565 7696 22664
rect 8036 22664 11376 22692
rect 11885 22695 11943 22701
rect 8036 22636 8064 22664
rect 11885 22661 11897 22695
rect 11931 22661 11943 22695
rect 11885 22655 11943 22661
rect 12342 22652 12348 22704
rect 12400 22652 12406 22704
rect 15654 22692 15660 22704
rect 14016 22664 15660 22692
rect 8018 22584 8024 22636
rect 8076 22584 8082 22636
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 8343 22596 8585 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 7653 22559 7711 22565
rect 7653 22525 7665 22559
rect 7699 22525 7711 22559
rect 7653 22519 7711 22525
rect 4430 22488 4436 22500
rect 3528 22460 4436 22488
rect 2961 22451 3019 22457
rect 4430 22448 4436 22460
rect 4488 22448 4494 22500
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 7101 22491 7159 22497
rect 7101 22457 7113 22491
rect 7147 22488 7159 22491
rect 8128 22488 8156 22587
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 11296 22596 11621 22624
rect 11296 22584 11302 22596
rect 11609 22593 11621 22596
rect 11655 22593 11667 22627
rect 11609 22587 11667 22593
rect 9674 22516 9680 22568
rect 9732 22556 9738 22568
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9732 22528 9781 22556
rect 9732 22516 9738 22528
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 9769 22519 9827 22525
rect 13630 22516 13636 22568
rect 13688 22516 13694 22568
rect 14016 22556 14044 22664
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22624 14151 22627
rect 14829 22627 14887 22633
rect 14139 22596 14780 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 14277 22559 14335 22565
rect 14277 22556 14289 22559
rect 14016 22528 14289 22556
rect 7147 22460 8156 22488
rect 7147 22457 7159 22460
rect 7101 22451 7159 22457
rect 934 22380 940 22432
rect 992 22420 998 22432
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 992 22392 1593 22420
rect 992 22380 998 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 2222 22380 2228 22432
rect 2280 22420 2286 22432
rect 2409 22423 2467 22429
rect 2409 22420 2421 22423
rect 2280 22392 2421 22420
rect 2280 22380 2286 22392
rect 2409 22389 2421 22392
rect 2455 22389 2467 22423
rect 2409 22383 2467 22389
rect 4522 22380 4528 22432
rect 4580 22380 4586 22432
rect 7024 22420 7052 22451
rect 8202 22448 8208 22500
rect 8260 22488 8266 22500
rect 8260 22460 9674 22488
rect 8260 22448 8266 22460
rect 8938 22420 8944 22432
rect 7024 22392 8944 22420
rect 8938 22380 8944 22392
rect 8996 22380 9002 22432
rect 9646 22420 9674 22460
rect 10134 22448 10140 22500
rect 10192 22448 10198 22500
rect 14108 22488 14136 22528
rect 14277 22525 14289 22528
rect 14323 22525 14335 22559
rect 14277 22519 14335 22525
rect 14550 22516 14556 22568
rect 14608 22556 14614 22568
rect 14645 22559 14703 22565
rect 14645 22556 14657 22559
rect 14608 22528 14657 22556
rect 14608 22516 14614 22528
rect 14645 22525 14657 22528
rect 14691 22525 14703 22559
rect 14752 22556 14780 22596
rect 14829 22593 14841 22627
rect 14875 22624 14887 22627
rect 15930 22624 15936 22636
rect 14875 22596 15936 22624
rect 14875 22593 14887 22596
rect 14829 22587 14887 22593
rect 15930 22584 15936 22596
rect 15988 22584 15994 22636
rect 15746 22556 15752 22568
rect 14752 22528 15752 22556
rect 14645 22519 14703 22525
rect 15746 22516 15752 22528
rect 15804 22556 15810 22568
rect 16040 22556 16068 22732
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 17460 22732 17785 22760
rect 17460 22720 17466 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 17773 22723 17831 22729
rect 19702 22720 19708 22772
rect 19760 22720 19766 22772
rect 21453 22763 21511 22769
rect 21453 22729 21465 22763
rect 21499 22760 21511 22763
rect 21910 22760 21916 22772
rect 21499 22732 21916 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 17494 22692 17500 22704
rect 16132 22664 17500 22692
rect 16132 22633 16160 22664
rect 17494 22652 17500 22664
rect 17552 22692 17558 22704
rect 17865 22695 17923 22701
rect 17865 22692 17877 22695
rect 17552 22664 17877 22692
rect 17552 22652 17558 22664
rect 17865 22661 17877 22664
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 16117 22627 16175 22633
rect 16117 22593 16129 22627
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 17770 22624 17776 22636
rect 16853 22587 16911 22593
rect 17236 22596 17776 22624
rect 15804 22528 16068 22556
rect 15804 22516 15810 22528
rect 16206 22516 16212 22568
rect 16264 22516 16270 22568
rect 16761 22559 16819 22565
rect 16761 22525 16773 22559
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 13556 22460 14136 22488
rect 13556 22420 13584 22460
rect 14182 22448 14188 22500
rect 14240 22488 14246 22500
rect 16485 22491 16543 22497
rect 16485 22488 16497 22491
rect 14240 22460 16497 22488
rect 14240 22448 14246 22460
rect 16485 22457 16497 22460
rect 16531 22457 16543 22491
rect 16485 22451 16543 22457
rect 9646 22392 13584 22420
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 16206 22420 16212 22432
rect 13688 22392 16212 22420
rect 13688 22380 13694 22392
rect 16206 22380 16212 22392
rect 16264 22420 16270 22432
rect 16776 22420 16804 22519
rect 16868 22488 16896 22587
rect 17236 22565 17264 22596
rect 17770 22584 17776 22596
rect 17828 22624 17834 22636
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 17828 22596 18061 22624
rect 17828 22584 17834 22596
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 19334 22584 19340 22636
rect 19392 22584 19398 22636
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 19720 22624 19748 22720
rect 20990 22652 20996 22704
rect 21048 22652 21054 22704
rect 19659 22596 19748 22624
rect 25501 22627 25559 22633
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 25501 22593 25513 22627
rect 25547 22593 25559 22627
rect 25501 22587 25559 22593
rect 17221 22559 17279 22565
rect 17221 22525 17233 22559
rect 17267 22525 17279 22559
rect 17221 22519 17279 22525
rect 17310 22516 17316 22568
rect 17368 22516 17374 22568
rect 17586 22516 17592 22568
rect 17644 22556 17650 22568
rect 18233 22559 18291 22565
rect 18233 22556 18245 22559
rect 17644 22528 18245 22556
rect 17644 22516 17650 22528
rect 18233 22525 18245 22528
rect 18279 22525 18291 22559
rect 19352 22556 19380 22584
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 19352 22528 19717 22556
rect 18233 22519 18291 22525
rect 19705 22525 19717 22528
rect 19751 22525 19763 22559
rect 19705 22519 19763 22525
rect 19981 22559 20039 22565
rect 19981 22525 19993 22559
rect 20027 22556 20039 22559
rect 20714 22556 20720 22568
rect 20027 22528 20720 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20714 22516 20720 22528
rect 20772 22516 20778 22568
rect 25516 22556 25544 22587
rect 25958 22556 25964 22568
rect 25516 22528 25964 22556
rect 25958 22516 25964 22528
rect 26016 22516 26022 22568
rect 17402 22488 17408 22500
rect 16868 22460 17408 22488
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 16264 22392 16804 22420
rect 16264 22380 16270 22392
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17604 22420 17632 22516
rect 17681 22491 17739 22497
rect 17681 22457 17693 22491
rect 17727 22457 17739 22491
rect 17681 22451 17739 22457
rect 17000 22392 17632 22420
rect 17696 22420 17724 22451
rect 18046 22420 18052 22432
rect 17696 22392 18052 22420
rect 17000 22380 17006 22392
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 19429 22423 19487 22429
rect 19429 22389 19441 22423
rect 19475 22420 19487 22423
rect 19978 22420 19984 22432
rect 19475 22392 19984 22420
rect 19475 22389 19487 22392
rect 19429 22383 19487 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 25317 22423 25375 22429
rect 25317 22389 25329 22423
rect 25363 22420 25375 22423
rect 26234 22420 26240 22432
rect 25363 22392 26240 22420
rect 25363 22389 25375 22392
rect 25317 22383 25375 22389
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 1104 22330 25852 22352
rect 1104 22278 4043 22330
rect 4095 22278 4107 22330
rect 4159 22278 4171 22330
rect 4223 22278 4235 22330
rect 4287 22278 4299 22330
rect 4351 22278 10230 22330
rect 10282 22278 10294 22330
rect 10346 22278 10358 22330
rect 10410 22278 10422 22330
rect 10474 22278 10486 22330
rect 10538 22278 16417 22330
rect 16469 22278 16481 22330
rect 16533 22278 16545 22330
rect 16597 22278 16609 22330
rect 16661 22278 16673 22330
rect 16725 22278 22604 22330
rect 22656 22278 22668 22330
rect 22720 22278 22732 22330
rect 22784 22278 22796 22330
rect 22848 22278 22860 22330
rect 22912 22278 25852 22330
rect 1104 22256 25852 22278
rect 2120 22219 2178 22225
rect 2120 22185 2132 22219
rect 2166 22216 2178 22219
rect 2222 22216 2228 22228
rect 2166 22188 2228 22216
rect 2166 22185 2178 22188
rect 2120 22179 2178 22185
rect 2222 22176 2228 22188
rect 2280 22176 2286 22228
rect 3602 22176 3608 22228
rect 3660 22176 3666 22228
rect 3786 22176 3792 22228
rect 3844 22176 3850 22228
rect 4430 22176 4436 22228
rect 4488 22176 4494 22228
rect 5445 22219 5503 22225
rect 5445 22185 5457 22219
rect 5491 22216 5503 22219
rect 5810 22216 5816 22228
rect 5491 22188 5816 22216
rect 5491 22185 5503 22188
rect 5445 22179 5503 22185
rect 5810 22176 5816 22188
rect 5868 22176 5874 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7101 22219 7159 22225
rect 7101 22216 7113 22219
rect 6972 22188 7113 22216
rect 6972 22176 6978 22188
rect 7101 22185 7113 22188
rect 7147 22185 7159 22219
rect 7101 22179 7159 22185
rect 7282 22176 7288 22228
rect 7340 22176 7346 22228
rect 7558 22176 7564 22228
rect 7616 22216 7622 22228
rect 10226 22216 10232 22228
rect 7616 22188 10232 22216
rect 7616 22176 7622 22188
rect 10226 22176 10232 22188
rect 10284 22176 10290 22228
rect 12250 22176 12256 22228
rect 12308 22176 12314 22228
rect 12342 22176 12348 22228
rect 12400 22176 12406 22228
rect 12894 22176 12900 22228
rect 12952 22216 12958 22228
rect 13630 22216 13636 22228
rect 12952 22188 13636 22216
rect 12952 22176 12958 22188
rect 13630 22176 13636 22188
rect 13688 22176 13694 22228
rect 14090 22176 14096 22228
rect 14148 22216 14154 22228
rect 14350 22219 14408 22225
rect 14350 22216 14362 22219
rect 14148 22188 14362 22216
rect 14148 22176 14154 22188
rect 14350 22185 14362 22188
rect 14396 22185 14408 22219
rect 14350 22179 14408 22185
rect 15930 22176 15936 22228
rect 15988 22176 15994 22228
rect 16298 22176 16304 22228
rect 16356 22216 16362 22228
rect 16356 22188 17264 22216
rect 16356 22176 16362 22188
rect 4448 22148 4476 22176
rect 5350 22148 5356 22160
rect 4448 22120 5356 22148
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4448 22080 4476 22120
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 7300 22148 7328 22176
rect 8662 22148 8668 22160
rect 6886 22120 7328 22148
rect 8496 22120 8668 22148
rect 4387 22052 4476 22080
rect 6457 22083 6515 22089
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 6457 22049 6469 22083
rect 6503 22080 6515 22083
rect 6886 22080 6914 22120
rect 6503 22052 6914 22080
rect 6503 22049 6515 22052
rect 6457 22043 6515 22049
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 21981 1915 22015
rect 1857 21975 1915 21981
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 22012 4767 22015
rect 5721 22015 5779 22021
rect 5721 22012 5733 22015
rect 4755 21984 5212 22012
rect 4755 21981 4767 21984
rect 4709 21975 4767 21981
rect 1872 21876 1900 21975
rect 5184 21956 5212 21984
rect 5644 21984 5733 22012
rect 2130 21904 2136 21956
rect 2188 21944 2194 21956
rect 4157 21947 4215 21953
rect 2188 21916 2622 21944
rect 2188 21904 2194 21916
rect 4157 21913 4169 21947
rect 4203 21944 4215 21947
rect 4430 21944 4436 21956
rect 4203 21916 4436 21944
rect 4203 21913 4215 21916
rect 4157 21907 4215 21913
rect 4430 21904 4436 21916
rect 4488 21904 4494 21956
rect 5166 21904 5172 21956
rect 5224 21904 5230 21956
rect 5644 21888 5672 21984
rect 5721 21981 5733 21984
rect 5767 21981 5779 22015
rect 5721 21975 5779 21981
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 6089 22015 6147 22021
rect 6089 22012 6101 22015
rect 5868 21984 6101 22012
rect 5868 21972 5874 21984
rect 6089 21981 6101 21984
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 2406 21876 2412 21888
rect 1872 21848 2412 21876
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 4249 21879 4307 21885
rect 4249 21845 4261 21879
rect 4295 21876 4307 21879
rect 5261 21879 5319 21885
rect 5261 21876 5273 21879
rect 4295 21848 5273 21876
rect 4295 21845 4307 21848
rect 4249 21839 4307 21845
rect 5261 21845 5273 21848
rect 5307 21845 5319 21879
rect 5261 21839 5319 21845
rect 5626 21836 5632 21888
rect 5684 21836 5690 21888
rect 5718 21836 5724 21888
rect 5776 21876 5782 21888
rect 5813 21879 5871 21885
rect 5813 21876 5825 21879
rect 5776 21848 5825 21876
rect 5776 21836 5782 21848
rect 5813 21845 5825 21848
rect 5859 21845 5871 21879
rect 5813 21839 5871 21845
rect 5902 21836 5908 21888
rect 5960 21836 5966 21888
rect 6196 21876 6224 21975
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 6696 21984 6776 22012
rect 6696 21972 6702 21984
rect 6748 21944 6776 21984
rect 6822 21972 6828 22024
rect 6880 22012 6886 22024
rect 7009 22015 7067 22021
rect 7009 22012 7021 22015
rect 6880 21984 7021 22012
rect 6880 21972 6886 21984
rect 7009 21981 7021 21984
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7116 21944 7144 21975
rect 7282 21972 7288 22024
rect 7340 21972 7346 22024
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 8496 22021 8524 22120
rect 8662 22108 8668 22120
rect 8720 22108 8726 22160
rect 9033 22151 9091 22157
rect 9033 22148 9045 22151
rect 8772 22120 9045 22148
rect 8772 22080 8800 22120
rect 9033 22117 9045 22120
rect 9079 22117 9091 22151
rect 9033 22111 9091 22117
rect 12069 22151 12127 22157
rect 12069 22117 12081 22151
rect 12115 22148 12127 22151
rect 12268 22148 12296 22176
rect 12989 22151 13047 22157
rect 12989 22148 13001 22151
rect 12115 22120 13001 22148
rect 12115 22117 12127 22120
rect 12069 22111 12127 22117
rect 12989 22117 13001 22120
rect 13035 22148 13047 22151
rect 13541 22151 13599 22157
rect 13541 22148 13553 22151
rect 13035 22120 13553 22148
rect 13035 22117 13047 22120
rect 12989 22111 13047 22117
rect 13541 22117 13553 22120
rect 13587 22117 13599 22151
rect 13541 22111 13599 22117
rect 15654 22108 15660 22160
rect 15712 22148 15718 22160
rect 15712 22120 16528 22148
rect 15712 22108 15718 22120
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 8588 22052 8800 22080
rect 8864 22052 9229 22080
rect 8588 22021 8616 22052
rect 8864 22024 8892 22052
rect 9217 22049 9229 22052
rect 9263 22049 9275 22083
rect 9217 22043 9275 22049
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 11606 22080 11612 22092
rect 10192 22052 11612 22080
rect 10192 22040 10198 22052
rect 11606 22040 11612 22052
rect 11664 22080 11670 22092
rect 12158 22080 12164 22092
rect 11664 22052 12164 22080
rect 11664 22040 11670 22052
rect 12158 22040 12164 22052
rect 12216 22040 12222 22092
rect 16500 22089 16528 22120
rect 12253 22083 12311 22089
rect 12253 22049 12265 22083
rect 12299 22080 12311 22083
rect 16485 22083 16543 22089
rect 12299 22052 12434 22080
rect 12299 22049 12311 22052
rect 12253 22043 12311 22049
rect 8389 22015 8447 22021
rect 8389 22012 8401 22015
rect 8352 21984 8401 22012
rect 8352 21972 8358 21984
rect 8389 21981 8401 21984
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 21981 8539 22015
rect 8481 21975 8539 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 8846 21972 8852 22024
rect 8904 21972 8910 22024
rect 8938 21972 8944 22024
rect 8996 21972 9002 22024
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 10778 21972 10784 22024
rect 10836 22012 10842 22024
rect 10836 21984 11284 22012
rect 10836 21972 10842 21984
rect 6748 21916 7144 21944
rect 8113 21947 8171 21953
rect 8113 21913 8125 21947
rect 8159 21944 8171 21947
rect 9493 21947 9551 21953
rect 9493 21944 9505 21947
rect 8159 21916 9505 21944
rect 8159 21913 8171 21916
rect 8113 21907 8171 21913
rect 9493 21913 9505 21916
rect 9539 21913 9551 21947
rect 10718 21916 11192 21944
rect 9493 21907 9551 21913
rect 6546 21876 6552 21888
rect 6196 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 6917 21879 6975 21885
rect 6917 21845 6929 21879
rect 6963 21876 6975 21879
rect 9582 21876 9588 21888
rect 6963 21848 9588 21876
rect 6963 21845 6975 21848
rect 6917 21839 6975 21845
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 10778 21836 10784 21888
rect 10836 21876 10842 21888
rect 11164 21885 11192 21916
rect 10965 21879 11023 21885
rect 10965 21876 10977 21879
rect 10836 21848 10977 21876
rect 10836 21836 10842 21848
rect 10965 21845 10977 21848
rect 11011 21845 11023 21879
rect 10965 21839 11023 21845
rect 11149 21879 11207 21885
rect 11149 21845 11161 21879
rect 11195 21845 11207 21879
rect 11256 21876 11284 21984
rect 11330 21972 11336 22024
rect 11388 21972 11394 22024
rect 11790 21972 11796 22024
rect 11848 21972 11854 22024
rect 12406 22012 12434 22052
rect 16485 22049 16497 22083
rect 16531 22080 16543 22083
rect 16531 22052 16565 22080
rect 16531 22049 16543 22052
rect 16485 22043 16543 22049
rect 17034 22040 17040 22092
rect 17092 22040 17098 22092
rect 17236 22080 17264 22188
rect 17310 22176 17316 22228
rect 17368 22216 17374 22228
rect 17678 22216 17684 22228
rect 17368 22188 17684 22216
rect 17368 22176 17374 22188
rect 17678 22176 17684 22188
rect 17736 22176 17742 22228
rect 17862 22176 17868 22228
rect 17920 22176 17926 22228
rect 18984 22188 20668 22216
rect 17681 22083 17739 22089
rect 17681 22080 17693 22083
rect 17236 22052 17693 22080
rect 17681 22049 17693 22052
rect 17727 22049 17739 22083
rect 17681 22043 17739 22049
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12406 21984 12541 22012
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13780 21984 14105 22012
rect 13780 21972 13786 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 16206 21972 16212 22024
rect 16264 22012 16270 22024
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 16264 21984 16313 22012
rect 16264 21972 16270 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16758 21972 16764 22024
rect 16816 21972 16822 22024
rect 16942 21972 16948 22024
rect 17000 21972 17006 22024
rect 17126 21972 17132 22024
rect 17184 21972 17190 22024
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 22012 17371 22015
rect 17402 22012 17408 22024
rect 17359 21984 17408 22012
rect 17359 21981 17371 21984
rect 17313 21975 17371 21981
rect 17402 21972 17408 21984
rect 17460 22012 17466 22024
rect 17586 22012 17592 22024
rect 17460 21984 17592 22012
rect 17460 21972 17466 21984
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 17770 21972 17776 22024
rect 17828 21972 17834 22024
rect 17880 22012 17908 22176
rect 18984 22089 19012 22188
rect 20640 22160 20668 22188
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 21085 22219 21143 22225
rect 21085 22216 21097 22219
rect 20772 22188 21097 22216
rect 20772 22176 20778 22188
rect 21085 22185 21097 22188
rect 21131 22185 21143 22219
rect 21085 22179 21143 22185
rect 20622 22108 20628 22160
rect 20680 22108 20686 22160
rect 18969 22083 19027 22089
rect 18969 22049 18981 22083
rect 19015 22049 19027 22083
rect 18969 22043 19027 22049
rect 19242 22040 19248 22092
rect 19300 22040 19306 22092
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 17880 21984 18705 22012
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 25501 22015 25559 22021
rect 25501 21981 25513 22015
rect 25547 21981 25559 22015
rect 25501 21975 25559 21981
rect 11422 21904 11428 21956
rect 11480 21944 11486 21956
rect 11808 21944 11836 21972
rect 12713 21947 12771 21953
rect 12713 21944 12725 21947
rect 11480 21916 12725 21944
rect 11480 21904 11486 21916
rect 12713 21913 12725 21916
rect 12759 21944 12771 21947
rect 13265 21947 13323 21953
rect 13265 21944 13277 21947
rect 12759 21916 13277 21944
rect 12759 21913 12771 21916
rect 12713 21907 12771 21913
rect 13265 21913 13277 21916
rect 13311 21913 13323 21947
rect 13265 21907 13323 21913
rect 13630 21904 13636 21956
rect 13688 21944 13694 21956
rect 16393 21947 16451 21953
rect 13688 21916 14858 21944
rect 13688 21904 13694 21916
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16439 21916 18184 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 13078 21876 13084 21888
rect 11256 21848 13084 21876
rect 11149 21839 11207 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13170 21836 13176 21888
rect 13228 21836 13234 21888
rect 13725 21879 13783 21885
rect 13725 21845 13737 21879
rect 13771 21876 13783 21879
rect 13814 21876 13820 21888
rect 13771 21848 13820 21876
rect 13771 21845 13783 21848
rect 13725 21839 13783 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14458 21836 14464 21888
rect 14516 21876 14522 21888
rect 15841 21879 15899 21885
rect 15841 21876 15853 21879
rect 14516 21848 15853 21876
rect 14516 21836 14522 21848
rect 15841 21845 15853 21848
rect 15887 21876 15899 21879
rect 16850 21876 16856 21888
rect 15887 21848 16856 21876
rect 15887 21845 15899 21848
rect 15841 21839 15899 21845
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 17494 21836 17500 21888
rect 17552 21836 17558 21888
rect 18156 21885 18184 21916
rect 19518 21904 19524 21956
rect 19576 21904 19582 21956
rect 19978 21904 19984 21956
rect 20036 21904 20042 21956
rect 25516 21944 25544 21975
rect 25958 21944 25964 21956
rect 25516 21916 25964 21944
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 18141 21879 18199 21885
rect 18141 21845 18153 21879
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 18322 21836 18328 21888
rect 18380 21836 18386 21888
rect 18785 21879 18843 21885
rect 18785 21845 18797 21879
rect 18831 21876 18843 21879
rect 18966 21876 18972 21888
rect 18831 21848 18972 21876
rect 18831 21845 18843 21848
rect 18785 21839 18843 21845
rect 18966 21836 18972 21848
rect 19024 21836 19030 21888
rect 20530 21836 20536 21888
rect 20588 21876 20594 21888
rect 20993 21879 21051 21885
rect 20993 21876 21005 21879
rect 20588 21848 21005 21876
rect 20588 21836 20594 21848
rect 20993 21845 21005 21848
rect 21039 21845 21051 21879
rect 20993 21839 21051 21845
rect 25317 21879 25375 21885
rect 25317 21845 25329 21879
rect 25363 21876 25375 21879
rect 25363 21848 25912 21876
rect 25363 21845 25375 21848
rect 25317 21839 25375 21845
rect 1104 21786 25852 21808
rect 1104 21734 4703 21786
rect 4755 21734 4767 21786
rect 4819 21734 4831 21786
rect 4883 21734 4895 21786
rect 4947 21734 4959 21786
rect 5011 21734 10890 21786
rect 10942 21734 10954 21786
rect 11006 21734 11018 21786
rect 11070 21734 11082 21786
rect 11134 21734 11146 21786
rect 11198 21734 17077 21786
rect 17129 21734 17141 21786
rect 17193 21734 17205 21786
rect 17257 21734 17269 21786
rect 17321 21734 17333 21786
rect 17385 21734 23264 21786
rect 23316 21734 23328 21786
rect 23380 21734 23392 21786
rect 23444 21734 23456 21786
rect 23508 21734 23520 21786
rect 23572 21734 25852 21786
rect 1104 21712 25852 21734
rect 2130 21632 2136 21684
rect 2188 21632 2194 21684
rect 2406 21632 2412 21684
rect 2464 21672 2470 21684
rect 8386 21672 8392 21684
rect 2464 21644 8392 21672
rect 2464 21632 2470 21644
rect 8386 21632 8392 21644
rect 8444 21672 8450 21684
rect 8846 21672 8852 21684
rect 8444 21644 8852 21672
rect 8444 21632 8450 21644
rect 8846 21632 8852 21644
rect 8904 21672 8910 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8904 21644 9137 21672
rect 8904 21632 8910 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 10505 21675 10563 21681
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 11330 21672 11336 21684
rect 10551 21644 11336 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 13170 21632 13176 21684
rect 13228 21632 13234 21684
rect 13265 21675 13323 21681
rect 13265 21641 13277 21675
rect 13311 21672 13323 21675
rect 13311 21644 14136 21672
rect 13311 21641 13323 21644
rect 13265 21635 13323 21641
rect 1489 21539 1547 21545
rect 1489 21505 1501 21539
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 1504 21400 1532 21499
rect 2314 21496 2320 21548
rect 2372 21496 2378 21548
rect 2424 21545 2452 21632
rect 3326 21564 3332 21616
rect 3384 21564 3390 21616
rect 4522 21564 4528 21616
rect 4580 21564 4586 21616
rect 4709 21607 4767 21613
rect 4709 21573 4721 21607
rect 4755 21604 4767 21607
rect 5626 21604 5632 21616
rect 4755 21576 5632 21604
rect 4755 21573 4767 21576
rect 4709 21567 4767 21573
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 5721 21607 5779 21613
rect 5721 21573 5733 21607
rect 5767 21604 5779 21607
rect 5994 21604 6000 21616
rect 5767 21576 6000 21604
rect 5767 21573 5779 21576
rect 5721 21567 5779 21573
rect 5994 21564 6000 21576
rect 6052 21564 6058 21616
rect 6362 21604 6368 21616
rect 6196 21576 6368 21604
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21505 2467 21539
rect 4540 21536 4568 21564
rect 2409 21499 2467 21505
rect 3896 21508 4568 21536
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21468 2743 21471
rect 3896 21468 3924 21508
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21536 4859 21539
rect 5258 21536 5264 21548
rect 4847 21508 5264 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 5258 21496 5264 21508
rect 5316 21536 5322 21548
rect 5905 21539 5963 21545
rect 5905 21536 5917 21539
rect 5316 21508 5917 21536
rect 5316 21496 5322 21508
rect 5905 21505 5917 21508
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 6086 21496 6092 21548
rect 6144 21496 6150 21548
rect 6196 21545 6224 21576
rect 6362 21564 6368 21576
rect 6420 21564 6426 21616
rect 6748 21576 7052 21604
rect 6181 21539 6239 21545
rect 6181 21505 6193 21539
rect 6227 21505 6239 21539
rect 6181 21499 6239 21505
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 2731 21440 3924 21468
rect 4157 21471 4215 21477
rect 2731 21437 2743 21440
rect 2685 21431 2743 21437
rect 4157 21437 4169 21471
rect 4203 21468 4215 21471
rect 5166 21468 5172 21480
rect 4203 21440 5172 21468
rect 4203 21437 4215 21440
rect 4157 21431 4215 21437
rect 5166 21428 5172 21440
rect 5224 21428 5230 21480
rect 5718 21428 5724 21480
rect 5776 21468 5782 21480
rect 6104 21468 6132 21496
rect 5776 21440 6132 21468
rect 5776 21428 5782 21440
rect 6638 21428 6644 21480
rect 6696 21428 6702 21480
rect 1504 21372 2544 21400
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1581 21335 1639 21341
rect 1581 21332 1593 21335
rect 992 21304 1593 21332
rect 992 21292 998 21304
rect 1581 21301 1593 21304
rect 1627 21301 1639 21335
rect 2516 21332 2544 21372
rect 5534 21360 5540 21412
rect 5592 21360 5598 21412
rect 5629 21403 5687 21409
rect 5629 21369 5641 21403
rect 5675 21400 5687 21403
rect 5810 21400 5816 21412
rect 5675 21372 5816 21400
rect 5675 21369 5687 21372
rect 5629 21363 5687 21369
rect 5810 21360 5816 21372
rect 5868 21360 5874 21412
rect 6748 21409 6776 21576
rect 7024 21545 7052 21576
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 7190 21564 7196 21616
rect 7248 21604 7254 21616
rect 7377 21607 7435 21613
rect 7377 21604 7389 21607
rect 7248 21576 7389 21604
rect 7248 21564 7254 21576
rect 7377 21573 7389 21576
rect 7423 21573 7435 21607
rect 7650 21604 7656 21616
rect 7377 21567 7435 21573
rect 7484 21576 7656 21604
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21536 6883 21539
rect 7009 21539 7067 21545
rect 6871 21508 6960 21536
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 6932 21468 6960 21508
rect 7009 21505 7021 21539
rect 7055 21505 7067 21539
rect 7116 21536 7144 21564
rect 7484 21545 7512 21576
rect 7650 21564 7656 21576
rect 7708 21564 7714 21616
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 10778 21604 10784 21616
rect 10008 21576 10784 21604
rect 10008 21564 10014 21576
rect 10778 21564 10784 21576
rect 10836 21564 10842 21616
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 7116 21508 7297 21536
rect 7009 21499 7067 21505
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7098 21468 7104 21480
rect 6932 21440 7104 21468
rect 7098 21428 7104 21440
rect 7156 21468 7162 21480
rect 7484 21468 7512 21499
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 12250 21536 12256 21548
rect 9640 21508 12256 21536
rect 9640 21496 9646 21508
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 13188 21536 13216 21632
rect 13722 21604 13728 21616
rect 13556 21576 13728 21604
rect 13556 21545 13584 21576
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 14108 21604 14136 21644
rect 16206 21632 16212 21684
rect 16264 21632 16270 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 17313 21675 17371 21681
rect 17313 21672 17325 21675
rect 16816 21644 17325 21672
rect 16816 21632 16822 21644
rect 17313 21641 17325 21644
rect 17359 21641 17371 21675
rect 17313 21635 17371 21641
rect 17865 21675 17923 21681
rect 17865 21641 17877 21675
rect 17911 21641 17923 21675
rect 17865 21635 17923 21641
rect 18601 21675 18659 21681
rect 18601 21641 18613 21675
rect 18647 21672 18659 21675
rect 19518 21672 19524 21684
rect 18647 21644 19524 21672
rect 18647 21641 18659 21644
rect 18601 21635 18659 21641
rect 14108 21576 14306 21604
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 13188 21508 13461 21536
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 13541 21539 13599 21545
rect 13541 21505 13553 21539
rect 13587 21505 13599 21539
rect 16224 21536 16252 21632
rect 16666 21564 16672 21616
rect 16724 21604 16730 21616
rect 17880 21604 17908 21635
rect 19518 21632 19524 21644
rect 19576 21632 19582 21684
rect 20073 21675 20131 21681
rect 20073 21641 20085 21675
rect 20119 21672 20131 21675
rect 21266 21672 21272 21684
rect 20119 21644 21272 21672
rect 20119 21641 20131 21644
rect 20073 21635 20131 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 23845 21675 23903 21681
rect 23845 21641 23857 21675
rect 23891 21672 23903 21675
rect 25884 21672 25912 21848
rect 23891 21644 25912 21672
rect 23891 21641 23903 21644
rect 23845 21635 23903 21641
rect 25222 21604 25228 21616
rect 16724 21576 17908 21604
rect 17972 21576 25228 21604
rect 16724 21564 16730 21576
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 16224 21508 16313 21536
rect 13541 21499 13599 21505
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 16393 21539 16451 21545
rect 16393 21505 16405 21539
rect 16439 21536 16451 21539
rect 16942 21536 16948 21548
rect 16439 21508 16948 21536
rect 16439 21505 16451 21508
rect 16393 21499 16451 21505
rect 16942 21496 16948 21508
rect 17000 21536 17006 21548
rect 17129 21539 17187 21545
rect 17129 21536 17141 21539
rect 17000 21508 17141 21536
rect 17000 21496 17006 21508
rect 17129 21505 17141 21508
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17972 21536 18000 21576
rect 25222 21564 25228 21576
rect 25280 21564 25286 21616
rect 17276 21508 18000 21536
rect 17276 21496 17282 21508
rect 18322 21496 18328 21548
rect 18380 21536 18386 21548
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18380 21508 18797 21536
rect 18380 21496 18386 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 20162 21496 20168 21548
rect 20220 21536 20226 21548
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 20220 21508 20453 21536
rect 20220 21496 20226 21508
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 21634 21496 21640 21548
rect 21692 21496 21698 21548
rect 21818 21496 21824 21548
rect 21876 21536 21882 21548
rect 21876 21508 24164 21536
rect 21876 21496 21882 21508
rect 24136 21480 24164 21508
rect 7156 21440 7512 21468
rect 7156 21428 7162 21440
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9732 21440 10057 21468
rect 9732 21428 9738 21440
rect 10045 21437 10057 21440
rect 10091 21437 10103 21471
rect 12802 21468 12808 21480
rect 10045 21431 10103 21437
rect 10152 21440 12808 21468
rect 6733 21403 6791 21409
rect 6733 21369 6745 21403
rect 6779 21369 6791 21403
rect 6733 21363 6791 21369
rect 4982 21332 4988 21344
rect 2516 21304 4988 21332
rect 1581 21295 1639 21301
rect 4982 21292 4988 21304
rect 5040 21292 5046 21344
rect 5828 21332 5856 21360
rect 6748 21332 6776 21363
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 10152 21400 10180 21440
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21468 13875 21471
rect 14182 21468 14188 21480
rect 13863 21440 14188 21468
rect 13863 21437 13875 21440
rect 13817 21431 13875 21437
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 17037 21471 17095 21477
rect 17037 21437 17049 21471
rect 17083 21437 17095 21471
rect 17037 21431 17095 21437
rect 7616 21372 10180 21400
rect 10321 21403 10379 21409
rect 7616 21360 7622 21372
rect 10321 21369 10333 21403
rect 10367 21369 10379 21403
rect 10321 21363 10379 21369
rect 15289 21403 15347 21409
rect 15289 21369 15301 21403
rect 15335 21400 15347 21403
rect 15470 21400 15476 21412
rect 15335 21372 15476 21400
rect 15335 21369 15347 21372
rect 15289 21363 15347 21369
rect 5828 21304 6776 21332
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10336 21332 10364 21363
rect 15470 21360 15476 21372
rect 15528 21400 15534 21412
rect 16942 21400 16948 21412
rect 15528 21372 16948 21400
rect 15528 21360 15534 21372
rect 16942 21360 16948 21372
rect 17000 21360 17006 21412
rect 17046 21400 17074 21431
rect 17402 21428 17408 21480
rect 17460 21468 17466 21480
rect 18046 21468 18052 21480
rect 17460 21440 18052 21468
rect 17460 21428 17466 21440
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 20530 21468 20536 21480
rect 19484 21440 20536 21468
rect 19484 21428 19490 21440
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 20622 21428 20628 21480
rect 20680 21428 20686 21480
rect 23937 21471 23995 21477
rect 23937 21468 23949 21471
rect 21376 21440 23949 21468
rect 17586 21400 17592 21412
rect 17046 21372 17592 21400
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 17678 21360 17684 21412
rect 17736 21360 17742 21412
rect 20254 21360 20260 21412
rect 20312 21400 20318 21412
rect 20640 21400 20668 21428
rect 20312 21372 20668 21400
rect 20312 21360 20318 21372
rect 10192 21304 10364 21332
rect 10192 21292 10198 21304
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 21376 21332 21404 21440
rect 23937 21437 23949 21440
rect 23983 21437 23995 21471
rect 23937 21431 23995 21437
rect 24118 21428 24124 21480
rect 24176 21428 24182 21480
rect 13136 21304 21404 21332
rect 13136 21292 13142 21304
rect 21450 21292 21456 21344
rect 21508 21292 21514 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23658 21332 23664 21344
rect 23523 21304 23664 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 1104 21242 25852 21264
rect 1104 21190 4043 21242
rect 4095 21190 4107 21242
rect 4159 21190 4171 21242
rect 4223 21190 4235 21242
rect 4287 21190 4299 21242
rect 4351 21190 10230 21242
rect 10282 21190 10294 21242
rect 10346 21190 10358 21242
rect 10410 21190 10422 21242
rect 10474 21190 10486 21242
rect 10538 21190 16417 21242
rect 16469 21190 16481 21242
rect 16533 21190 16545 21242
rect 16597 21190 16609 21242
rect 16661 21190 16673 21242
rect 16725 21190 22604 21242
rect 22656 21190 22668 21242
rect 22720 21190 22732 21242
rect 22784 21190 22796 21242
rect 22848 21190 22860 21242
rect 22912 21190 25852 21242
rect 1104 21168 25852 21190
rect 2314 21088 2320 21140
rect 2372 21128 2378 21140
rect 2685 21131 2743 21137
rect 2685 21128 2697 21131
rect 2372 21100 2697 21128
rect 2372 21088 2378 21100
rect 2685 21097 2697 21100
rect 2731 21097 2743 21131
rect 2685 21091 2743 21097
rect 3234 21088 3240 21140
rect 3292 21088 3298 21140
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 5445 21131 5503 21137
rect 5445 21097 5457 21131
rect 5491 21128 5503 21131
rect 5534 21128 5540 21140
rect 5491 21100 5540 21128
rect 5491 21097 5503 21100
rect 5445 21091 5503 21097
rect 5534 21088 5540 21100
rect 5592 21088 5598 21140
rect 6546 21088 6552 21140
rect 6604 21128 6610 21140
rect 7282 21128 7288 21140
rect 6604 21100 7288 21128
rect 6604 21088 6610 21100
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 11241 21131 11299 21137
rect 9646 21100 10640 21128
rect 2593 21063 2651 21069
rect 2593 21029 2605 21063
rect 2639 21060 2651 21063
rect 3145 21063 3203 21069
rect 3145 21060 3157 21063
rect 2639 21032 3157 21060
rect 2639 21029 2651 21032
rect 2593 21023 2651 21029
rect 3145 21029 3157 21032
rect 3191 21060 3203 21063
rect 3252 21060 3280 21088
rect 3191 21032 3280 21060
rect 5629 21063 5687 21069
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 5629 21029 5641 21063
rect 5675 21060 5687 21063
rect 5902 21060 5908 21072
rect 5675 21032 5908 21060
rect 5675 21029 5687 21032
rect 5629 21023 5687 21029
rect 5902 21020 5908 21032
rect 5960 21060 5966 21072
rect 7098 21060 7104 21072
rect 5960 21032 7104 21060
rect 5960 21020 5966 21032
rect 7098 21020 7104 21032
rect 7156 21020 7162 21072
rect 9646 21060 9674 21100
rect 7208 21032 9674 21060
rect 10045 21063 10103 21069
rect 3237 20995 3295 21001
rect 3237 20961 3249 20995
rect 3283 20961 3295 20995
rect 3237 20955 3295 20961
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 3252 20924 3280 20955
rect 4430 20952 4436 21004
rect 4488 20992 4494 21004
rect 7208 20992 7236 21032
rect 10045 21029 10057 21063
rect 10091 21060 10103 21063
rect 10134 21060 10140 21072
rect 10091 21032 10140 21060
rect 10091 21029 10103 21032
rect 10045 21023 10103 21029
rect 10134 21020 10140 21032
rect 10192 21060 10198 21072
rect 10505 21063 10563 21069
rect 10505 21060 10517 21063
rect 10192 21032 10517 21060
rect 10192 21020 10198 21032
rect 10505 21029 10517 21032
rect 10551 21029 10563 21063
rect 10612 21060 10640 21100
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11422 21128 11428 21140
rect 11287 21100 11428 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 11422 21088 11428 21100
rect 11480 21088 11486 21140
rect 11606 21088 11612 21140
rect 11664 21088 11670 21140
rect 11716 21100 12434 21128
rect 11716 21060 11744 21100
rect 10612 21032 11744 21060
rect 10505 21023 10563 21029
rect 11790 21020 11796 21072
rect 11848 21060 11854 21072
rect 12161 21063 12219 21069
rect 12161 21060 12173 21063
rect 11848 21032 12173 21060
rect 11848 21020 11854 21032
rect 12161 21029 12173 21032
rect 12207 21029 12219 21063
rect 12406 21060 12434 21100
rect 13630 21088 13636 21140
rect 13688 21088 13694 21140
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 17129 21131 17187 21137
rect 17129 21128 17141 21131
rect 13780 21100 17141 21128
rect 13780 21088 13786 21100
rect 17129 21097 17141 21100
rect 17175 21128 17187 21131
rect 19334 21128 19340 21140
rect 17175 21100 19340 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 20809 21131 20867 21137
rect 20809 21097 20821 21131
rect 20855 21128 20867 21131
rect 21634 21128 21640 21140
rect 20855 21100 21640 21128
rect 20855 21097 20867 21100
rect 20809 21091 20867 21097
rect 21634 21088 21640 21100
rect 21692 21088 21698 21140
rect 12406 21032 17264 21060
rect 12161 21023 12219 21029
rect 4488 20964 7236 20992
rect 4488 20952 4494 20964
rect 7834 20952 7840 21004
rect 7892 20992 7898 21004
rect 17236 20992 17264 21032
rect 20622 21020 20628 21072
rect 20680 21020 20686 21072
rect 25501 21063 25559 21069
rect 25501 21029 25513 21063
rect 25547 21060 25559 21063
rect 26326 21060 26332 21072
rect 25547 21032 26332 21060
rect 25547 21029 25559 21032
rect 25501 21023 25559 21029
rect 26326 21020 26332 21032
rect 26384 21020 26390 21072
rect 24946 20992 24952 21004
rect 7892 20964 15700 20992
rect 17236 20964 24952 20992
rect 7892 20952 7898 20964
rect 3513 20927 3571 20933
rect 3513 20924 3525 20927
rect 3252 20896 3525 20924
rect 3513 20893 3525 20896
rect 3559 20893 3571 20927
rect 3513 20887 3571 20893
rect 5166 20884 5172 20936
rect 5224 20884 5230 20936
rect 5258 20884 5264 20936
rect 5316 20924 5322 20936
rect 5534 20924 5540 20936
rect 5316 20896 5540 20924
rect 5316 20884 5322 20896
rect 5534 20884 5540 20896
rect 5592 20924 5598 20936
rect 8294 20924 8300 20936
rect 5592 20896 8300 20924
rect 5592 20884 5598 20896
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20893 8815 20927
rect 8757 20887 8815 20893
rect 2225 20859 2283 20865
rect 2225 20825 2237 20859
rect 2271 20856 2283 20859
rect 2777 20859 2835 20865
rect 2777 20856 2789 20859
rect 2271 20828 2789 20856
rect 2271 20825 2283 20828
rect 2225 20819 2283 20825
rect 2777 20825 2789 20828
rect 2823 20856 2835 20859
rect 2958 20856 2964 20868
rect 2823 20828 2964 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2958 20816 2964 20828
rect 3016 20816 3022 20868
rect 4982 20816 4988 20868
rect 5040 20856 5046 20868
rect 7558 20856 7564 20868
rect 5040 20828 7564 20856
rect 5040 20816 5046 20828
rect 7558 20816 7564 20828
rect 7616 20816 7622 20868
rect 8772 20856 8800 20887
rect 8938 20884 8944 20936
rect 8996 20884 9002 20936
rect 10318 20924 10324 20936
rect 9048 20896 10324 20924
rect 9048 20856 9076 20896
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 11422 20924 11428 20936
rect 10428 20896 11428 20924
rect 8772 20828 9076 20856
rect 9674 20816 9680 20868
rect 9732 20856 9738 20868
rect 10229 20859 10287 20865
rect 10229 20856 10241 20859
rect 9732 20828 10241 20856
rect 9732 20816 9738 20828
rect 10229 20825 10241 20828
rect 10275 20856 10287 20859
rect 10428 20856 10456 20896
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 13814 20884 13820 20936
rect 13872 20884 13878 20936
rect 14182 20884 14188 20936
rect 14240 20884 14246 20936
rect 14366 20884 14372 20936
rect 14424 20884 14430 20936
rect 14458 20884 14464 20936
rect 14516 20884 14522 20936
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 10275 20828 10456 20856
rect 11149 20859 11207 20865
rect 10275 20825 10287 20828
rect 10229 20819 10287 20825
rect 11149 20825 11161 20859
rect 11195 20856 11207 20859
rect 11238 20856 11244 20868
rect 11195 20828 11244 20856
rect 11195 20825 11207 20828
rect 11149 20819 11207 20825
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11514 20816 11520 20868
rect 11572 20816 11578 20868
rect 11882 20816 11888 20868
rect 11940 20856 11946 20868
rect 13170 20856 13176 20868
rect 11940 20828 13176 20856
rect 11940 20816 11946 20828
rect 13170 20816 13176 20828
rect 13228 20816 13234 20868
rect 1578 20748 1584 20800
rect 1636 20748 1642 20800
rect 6638 20748 6644 20800
rect 6696 20788 6702 20800
rect 7374 20788 7380 20800
rect 6696 20760 7380 20788
rect 6696 20748 6702 20760
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 8570 20748 8576 20800
rect 8628 20748 8634 20800
rect 9582 20748 9588 20800
rect 9640 20748 9646 20800
rect 10134 20748 10140 20800
rect 10192 20748 10198 20800
rect 10318 20748 10324 20800
rect 10376 20788 10382 20800
rect 10689 20791 10747 20797
rect 10689 20788 10701 20791
rect 10376 20760 10701 20788
rect 10376 20748 10382 20760
rect 10689 20757 10701 20760
rect 10735 20757 10747 20791
rect 10689 20751 10747 20757
rect 12345 20791 12403 20797
rect 12345 20757 12357 20791
rect 12391 20788 12403 20791
rect 12986 20788 12992 20800
rect 12391 20760 12992 20788
rect 12391 20757 12403 20760
rect 12345 20751 12403 20757
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 14200 20797 14228 20884
rect 14384 20856 14412 20884
rect 14568 20856 14596 20887
rect 14642 20884 14648 20936
rect 14700 20884 14706 20936
rect 14734 20884 14740 20936
rect 14792 20924 14798 20936
rect 15672 20933 15700 20964
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 14829 20927 14887 20933
rect 14829 20924 14841 20927
rect 14792 20896 14841 20924
rect 14792 20884 14798 20896
rect 14829 20893 14841 20896
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20924 15715 20927
rect 16206 20924 16212 20936
rect 15703 20896 16212 20924
rect 15703 20893 15715 20896
rect 15657 20887 15715 20893
rect 16206 20884 16212 20896
rect 16264 20884 16270 20936
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 20588 20896 20913 20924
rect 20588 20884 20594 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 25363 20896 26004 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 14384 20828 14596 20856
rect 14185 20791 14243 20797
rect 14185 20757 14197 20791
rect 14231 20757 14243 20791
rect 14185 20751 14243 20757
rect 14274 20748 14280 20800
rect 14332 20788 14338 20800
rect 14752 20788 14780 20884
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 20349 20859 20407 20865
rect 20349 20856 20361 20859
rect 19392 20828 20361 20856
rect 19392 20816 19398 20828
rect 20349 20825 20361 20828
rect 20395 20825 20407 20859
rect 20349 20819 20407 20825
rect 21174 20816 21180 20868
rect 21232 20816 21238 20868
rect 21450 20816 21456 20868
rect 21508 20856 21514 20868
rect 21508 20828 21666 20856
rect 21508 20816 21514 20828
rect 14332 20760 14780 20788
rect 14332 20748 14338 20760
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 22186 20788 22192 20800
rect 17460 20760 22192 20788
rect 17460 20748 17466 20760
rect 22186 20748 22192 20760
rect 22244 20788 22250 20800
rect 22649 20791 22707 20797
rect 22649 20788 22661 20791
rect 22244 20760 22661 20788
rect 22244 20748 22250 20760
rect 22649 20757 22661 20760
rect 22695 20757 22707 20791
rect 22649 20751 22707 20757
rect 25976 20732 26004 20896
rect 1104 20698 25852 20720
rect 1104 20646 4703 20698
rect 4755 20646 4767 20698
rect 4819 20646 4831 20698
rect 4883 20646 4895 20698
rect 4947 20646 4959 20698
rect 5011 20646 10890 20698
rect 10942 20646 10954 20698
rect 11006 20646 11018 20698
rect 11070 20646 11082 20698
rect 11134 20646 11146 20698
rect 11198 20646 17077 20698
rect 17129 20646 17141 20698
rect 17193 20646 17205 20698
rect 17257 20646 17269 20698
rect 17321 20646 17333 20698
rect 17385 20646 23264 20698
rect 23316 20646 23328 20698
rect 23380 20646 23392 20698
rect 23444 20646 23456 20698
rect 23508 20646 23520 20698
rect 23572 20646 25852 20698
rect 25958 20680 25964 20732
rect 26016 20680 26022 20732
rect 1104 20624 25852 20646
rect 2869 20587 2927 20593
rect 2869 20553 2881 20587
rect 2915 20584 2927 20587
rect 4798 20584 4804 20596
rect 2915 20556 4804 20584
rect 2915 20553 2927 20556
rect 2869 20547 2927 20553
rect 4798 20544 4804 20556
rect 4856 20544 4862 20596
rect 9582 20584 9588 20596
rect 7576 20556 9588 20584
rect 3234 20476 3240 20528
rect 3292 20516 3298 20528
rect 7576 20516 7604 20556
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 10134 20544 10140 20596
rect 10192 20544 10198 20596
rect 11241 20587 11299 20593
rect 11241 20553 11253 20587
rect 11287 20584 11299 20587
rect 11882 20584 11888 20596
rect 11287 20556 11888 20584
rect 11287 20553 11299 20556
rect 11241 20547 11299 20553
rect 9950 20516 9956 20528
rect 3292 20488 4108 20516
rect 3292 20476 3298 20488
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20380 2467 20383
rect 2958 20380 2964 20392
rect 2455 20352 2964 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 3712 20380 3740 20411
rect 3786 20408 3792 20460
rect 3844 20448 3850 20460
rect 3973 20451 4031 20457
rect 3973 20448 3985 20451
rect 3844 20420 3985 20448
rect 3844 20408 3850 20420
rect 3973 20417 3985 20420
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 3467 20352 3740 20380
rect 4080 20380 4108 20488
rect 7484 20488 7604 20516
rect 9890 20488 9956 20516
rect 7484 20457 7512 20488
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 7098 20380 7104 20392
rect 4080 20352 7104 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 7098 20340 7104 20352
rect 7156 20340 7162 20392
rect 7576 20380 7604 20411
rect 7650 20408 7656 20460
rect 7708 20408 7714 20460
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 8386 20408 8392 20460
rect 8444 20408 8450 20460
rect 10152 20448 10180 20544
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10152 20420 10517 20448
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 11057 20451 11115 20457
rect 11057 20417 11069 20451
rect 11103 20448 11115 20451
rect 11146 20448 11152 20460
rect 11103 20420 11152 20448
rect 11103 20417 11115 20420
rect 11057 20411 11115 20417
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 8662 20380 8668 20392
rect 7576 20352 8668 20380
rect 8662 20340 8668 20352
rect 8720 20380 8726 20392
rect 9306 20380 9312 20392
rect 8720 20352 9312 20380
rect 8720 20340 8726 20352
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 11256 20380 11284 20547
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12345 20587 12403 20593
rect 12345 20553 12357 20587
rect 12391 20584 12403 20587
rect 12710 20584 12716 20596
rect 12391 20556 12716 20584
rect 12391 20553 12403 20556
rect 12345 20547 12403 20553
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12802 20544 12808 20596
rect 12860 20544 12866 20596
rect 13170 20544 13176 20596
rect 13228 20544 13234 20596
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 21232 20556 21373 20584
rect 21232 20544 21238 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 21821 20587 21879 20593
rect 21821 20553 21833 20587
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 11514 20408 11520 20460
rect 11572 20448 11578 20460
rect 11882 20448 11888 20460
rect 11572 20420 11888 20448
rect 11572 20408 11578 20420
rect 11882 20408 11888 20420
rect 11940 20408 11946 20460
rect 12986 20408 12992 20460
rect 13044 20408 13050 20460
rect 13188 20448 13216 20544
rect 15841 20519 15899 20525
rect 15841 20485 15853 20519
rect 15887 20516 15899 20519
rect 16114 20516 16120 20528
rect 15887 20488 16120 20516
rect 15887 20485 15899 20488
rect 15841 20479 15899 20485
rect 16114 20476 16120 20488
rect 16172 20476 16178 20528
rect 13188 20420 15884 20448
rect 9692 20352 11284 20380
rect 12437 20383 12495 20389
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20312 2835 20315
rect 3234 20312 3240 20324
rect 2823 20284 3240 20312
rect 2823 20281 2835 20284
rect 2777 20275 2835 20281
rect 3234 20272 3240 20284
rect 3292 20272 3298 20324
rect 3510 20204 3516 20256
rect 3568 20204 3574 20256
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 3789 20247 3847 20253
rect 3789 20244 3801 20247
rect 3660 20216 3801 20244
rect 3660 20204 3666 20216
rect 3789 20213 3801 20216
rect 3835 20213 3847 20247
rect 3789 20207 3847 20213
rect 7190 20204 7196 20256
rect 7248 20204 7254 20256
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 8646 20247 8704 20253
rect 8646 20244 8658 20247
rect 8444 20216 8658 20244
rect 8444 20204 8450 20216
rect 8646 20213 8658 20216
rect 8692 20213 8704 20247
rect 8646 20207 8704 20213
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 9692 20244 9720 20352
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 15856 20380 15884 20420
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15988 20420 16037 20448
rect 15988 20408 15994 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16298 20448 16304 20460
rect 16255 20420 16304 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 20349 20451 20407 20457
rect 18463 20420 19334 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 18322 20380 18328 20392
rect 15856 20352 18328 20380
rect 18322 20340 18328 20352
rect 18380 20340 18386 20392
rect 19306 20380 19334 20420
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 20438 20448 20444 20460
rect 20395 20420 20444 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 21545 20451 21603 20457
rect 21545 20417 21557 20451
rect 21591 20448 21603 20451
rect 21836 20448 21864 20547
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 22281 20587 22339 20593
rect 22281 20584 22293 20587
rect 22244 20556 22293 20584
rect 22244 20544 22250 20556
rect 22281 20553 22293 20556
rect 22327 20553 22339 20587
rect 22281 20547 22339 20553
rect 23658 20544 23664 20596
rect 23716 20544 23722 20596
rect 21591 20420 21864 20448
rect 22189 20451 22247 20457
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22462 20448 22468 20460
rect 22235 20420 22468 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 22462 20408 22468 20420
rect 22520 20448 22526 20460
rect 23106 20448 23112 20460
rect 22520 20420 23112 20448
rect 22520 20408 22526 20420
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23676 20448 23704 20544
rect 23753 20451 23811 20457
rect 23753 20448 23765 20451
rect 23676 20420 23765 20448
rect 23753 20417 23765 20420
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 19794 20380 19800 20392
rect 19306 20352 19800 20380
rect 19794 20340 19800 20352
rect 19852 20380 19858 20392
rect 19852 20352 22094 20380
rect 19852 20340 19858 20352
rect 9950 20272 9956 20324
rect 10008 20312 10014 20324
rect 10321 20315 10379 20321
rect 10321 20312 10333 20315
rect 10008 20284 10333 20312
rect 10008 20272 10014 20284
rect 10321 20281 10333 20284
rect 10367 20281 10379 20315
rect 10321 20275 10379 20281
rect 11422 20272 11428 20324
rect 11480 20312 11486 20324
rect 11977 20315 12035 20321
rect 11977 20312 11989 20315
rect 11480 20284 11989 20312
rect 11480 20272 11486 20284
rect 11977 20281 11989 20284
rect 12023 20281 12035 20315
rect 11977 20275 12035 20281
rect 12250 20272 12256 20324
rect 12308 20312 12314 20324
rect 15378 20312 15384 20324
rect 12308 20284 15384 20312
rect 12308 20272 12314 20284
rect 15378 20272 15384 20284
rect 15436 20312 15442 20324
rect 15930 20312 15936 20324
rect 15436 20284 15936 20312
rect 15436 20272 15442 20284
rect 15930 20272 15936 20284
rect 15988 20272 15994 20324
rect 8904 20216 9720 20244
rect 8904 20204 8910 20216
rect 10134 20204 10140 20256
rect 10192 20204 10198 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 11698 20244 11704 20256
rect 11388 20216 11704 20244
rect 11388 20204 11394 20216
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 18598 20244 18604 20256
rect 12492 20216 18604 20244
rect 12492 20204 12498 20216
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 20128 20216 20545 20244
rect 20128 20204 20134 20216
rect 20533 20213 20545 20216
rect 20579 20213 20591 20247
rect 22066 20244 22094 20352
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 22186 20244 22192 20256
rect 22066 20216 22192 20244
rect 20533 20207 20591 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 23569 20247 23627 20253
rect 23569 20213 23581 20247
rect 23615 20244 23627 20247
rect 23658 20244 23664 20256
rect 23615 20216 23664 20244
rect 23615 20213 23627 20216
rect 23569 20207 23627 20213
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 1104 20154 25852 20176
rect 1104 20102 4043 20154
rect 4095 20102 4107 20154
rect 4159 20102 4171 20154
rect 4223 20102 4235 20154
rect 4287 20102 4299 20154
rect 4351 20102 10230 20154
rect 10282 20102 10294 20154
rect 10346 20102 10358 20154
rect 10410 20102 10422 20154
rect 10474 20102 10486 20154
rect 10538 20102 16417 20154
rect 16469 20102 16481 20154
rect 16533 20102 16545 20154
rect 16597 20102 16609 20154
rect 16661 20102 16673 20154
rect 16725 20102 22604 20154
rect 22656 20102 22668 20154
rect 22720 20102 22732 20154
rect 22784 20102 22796 20154
rect 22848 20102 22860 20154
rect 22912 20102 25852 20154
rect 1104 20080 25852 20102
rect 2590 20000 2596 20052
rect 2648 20040 2654 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 2648 20012 3801 20040
rect 2648 20000 2654 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 4062 20000 4068 20052
rect 4120 20040 4126 20052
rect 4617 20043 4675 20049
rect 4617 20040 4629 20043
rect 4120 20012 4629 20040
rect 4120 20000 4126 20012
rect 4617 20009 4629 20012
rect 4663 20009 4675 20043
rect 4617 20003 4675 20009
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 4764 20012 6316 20040
rect 4764 20000 4770 20012
rect 6288 19981 6316 20012
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 7009 20043 7067 20049
rect 7009 20040 7021 20043
rect 6696 20012 7021 20040
rect 6696 20000 6702 20012
rect 7009 20009 7021 20012
rect 7055 20040 7067 20043
rect 7282 20040 7288 20052
rect 7055 20012 7288 20040
rect 7055 20009 7067 20012
rect 7009 20003 7067 20009
rect 7282 20000 7288 20012
rect 7340 20000 7346 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 7745 20043 7803 20049
rect 7745 20040 7757 20043
rect 7708 20012 7757 20040
rect 7708 20000 7714 20012
rect 7745 20009 7757 20012
rect 7791 20009 7803 20043
rect 7745 20003 7803 20009
rect 8386 20000 8392 20052
rect 8444 20040 8450 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8444 20012 8953 20040
rect 8444 20000 8450 20012
rect 8941 20009 8953 20012
rect 8987 20009 8999 20043
rect 8941 20003 8999 20009
rect 9030 20000 9036 20052
rect 9088 20040 9094 20052
rect 9214 20040 9220 20052
rect 9088 20012 9220 20040
rect 9088 20000 9094 20012
rect 9214 20000 9220 20012
rect 9272 20040 9278 20052
rect 9674 20040 9680 20052
rect 9272 20012 9680 20040
rect 9272 20000 9278 20012
rect 9674 20000 9680 20012
rect 9732 20040 9738 20052
rect 10134 20040 10140 20052
rect 9732 20012 10140 20040
rect 9732 20000 9738 20012
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 11514 20040 11520 20052
rect 11204 20012 11520 20040
rect 11204 20000 11210 20012
rect 11514 20000 11520 20012
rect 11572 20040 11578 20052
rect 12434 20040 12440 20052
rect 11572 20012 12440 20040
rect 11572 20000 11578 20012
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 12584 20012 13277 20040
rect 12584 20000 12590 20012
rect 13265 20009 13277 20012
rect 13311 20040 13323 20043
rect 14182 20040 14188 20052
rect 13311 20012 14188 20040
rect 13311 20009 13323 20012
rect 13265 20003 13323 20009
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14700 20012 15025 20040
rect 14700 20000 14706 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15378 20000 15384 20052
rect 15436 20000 15442 20052
rect 16298 20040 16304 20052
rect 15580 20012 16304 20040
rect 5169 19975 5227 19981
rect 5169 19972 5181 19975
rect 3160 19944 5181 19972
rect 1670 19864 1676 19916
rect 1728 19904 1734 19916
rect 1765 19907 1823 19913
rect 1765 19904 1777 19907
rect 1728 19876 1777 19904
rect 1728 19864 1734 19876
rect 1765 19873 1777 19876
rect 1811 19904 1823 19907
rect 2682 19904 2688 19916
rect 1811 19876 2688 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 3160 19822 3188 19944
rect 5169 19941 5181 19944
rect 5215 19941 5227 19975
rect 5169 19935 5227 19941
rect 6273 19975 6331 19981
rect 6273 19941 6285 19975
rect 6319 19941 6331 19975
rect 6273 19935 6331 19941
rect 3694 19864 3700 19916
rect 3752 19904 3758 19916
rect 4062 19904 4068 19916
rect 3752 19876 4068 19904
rect 3752 19864 3758 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4246 19864 4252 19916
rect 4304 19904 4310 19916
rect 4341 19907 4399 19913
rect 4341 19904 4353 19907
rect 4304 19876 4353 19904
rect 4304 19864 4310 19876
rect 4341 19873 4353 19876
rect 4387 19873 4399 19907
rect 4341 19867 4399 19873
rect 4448 19904 4568 19912
rect 4709 19907 4767 19913
rect 4709 19904 4721 19907
rect 4448 19884 4721 19904
rect 4448 19848 4476 19884
rect 4540 19876 4721 19884
rect 4709 19873 4721 19876
rect 4755 19873 4767 19907
rect 4709 19867 4767 19873
rect 4798 19864 4804 19916
rect 4856 19904 4862 19916
rect 6288 19904 6316 19935
rect 6822 19932 6828 19984
rect 6880 19932 6886 19984
rect 7098 19932 7104 19984
rect 7156 19972 7162 19984
rect 11330 19972 11336 19984
rect 7156 19944 11336 19972
rect 7156 19932 7162 19944
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 4856 19876 5396 19904
rect 6288 19876 6561 19904
rect 4856 19864 4862 19876
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4203 19808 4384 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4356 19780 4384 19808
rect 4430 19796 4436 19848
rect 4488 19796 4494 19848
rect 4522 19796 4528 19848
rect 4580 19836 4586 19848
rect 4617 19839 4675 19845
rect 4617 19836 4629 19839
rect 4580 19808 4629 19836
rect 4580 19796 4586 19808
rect 4617 19805 4629 19808
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 5074 19836 5080 19848
rect 4893 19799 4951 19805
rect 5000 19808 5080 19836
rect 2038 19728 2044 19780
rect 2096 19728 2102 19780
rect 3528 19740 4292 19768
rect 3528 19709 3556 19740
rect 4264 19709 4292 19740
rect 4338 19728 4344 19780
rect 4396 19768 4402 19780
rect 4908 19768 4936 19799
rect 4396 19740 4936 19768
rect 4396 19728 4402 19740
rect 3513 19703 3571 19709
rect 3513 19669 3525 19703
rect 3559 19669 3571 19703
rect 3513 19663 3571 19669
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 5000 19700 5028 19808
rect 5074 19796 5080 19808
rect 5132 19796 5138 19848
rect 5368 19845 5396 19876
rect 6549 19873 6561 19876
rect 6595 19873 6607 19907
rect 6549 19867 6607 19873
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19836 6055 19839
rect 6840 19836 6868 19932
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 7760 19876 7849 19904
rect 6043 19808 6868 19836
rect 6043 19805 6055 19808
rect 5997 19799 6055 19805
rect 7098 19796 7104 19848
rect 7156 19796 7162 19848
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 6822 19728 6828 19780
rect 6880 19768 6886 19780
rect 7300 19768 7328 19799
rect 7374 19796 7380 19848
rect 7432 19836 7438 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 7432 19808 7481 19836
rect 7432 19796 7438 19808
rect 7469 19805 7481 19808
rect 7515 19836 7527 19839
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 7515 19808 7573 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 7650 19796 7656 19848
rect 7708 19796 7714 19848
rect 6880 19740 7328 19768
rect 6880 19728 6886 19740
rect 4295 19672 5028 19700
rect 5077 19703 5135 19709
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5442 19700 5448 19712
rect 5123 19672 5448 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 6454 19660 6460 19712
rect 6512 19660 6518 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7760 19700 7788 19876
rect 7837 19873 7849 19876
rect 7883 19873 7895 19907
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 7837 19867 7895 19873
rect 9048 19876 9628 19904
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19836 8539 19839
rect 8662 19836 8668 19848
rect 8527 19808 8668 19836
rect 8527 19805 8539 19808
rect 8481 19799 8539 19805
rect 7340 19672 7788 19700
rect 8312 19700 8340 19799
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 8754 19796 8760 19848
rect 8812 19836 8818 19848
rect 9048 19836 9076 19876
rect 8812 19808 9076 19836
rect 8812 19796 8818 19808
rect 9214 19796 9220 19848
rect 9272 19796 9278 19848
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9600 19845 9628 19876
rect 11348 19876 11529 19904
rect 11348 19848 11376 19876
rect 11517 19873 11529 19876
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 12526 19904 12532 19916
rect 11940 19876 12532 19904
rect 11940 19864 11946 19876
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 15102 19864 15108 19916
rect 15160 19864 15166 19916
rect 15396 19904 15424 20000
rect 15580 19904 15608 20012
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 17494 20040 17500 20052
rect 16807 20012 17500 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 15657 19975 15715 19981
rect 15657 19941 15669 19975
rect 15703 19972 15715 19975
rect 16114 19972 16120 19984
rect 15703 19944 16120 19972
rect 15703 19941 15715 19944
rect 15657 19935 15715 19941
rect 16114 19932 16120 19944
rect 16172 19932 16178 19984
rect 16776 19972 16804 20003
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18322 20000 18328 20052
rect 18380 20000 18386 20052
rect 25409 20043 25467 20049
rect 25409 20009 25421 20043
rect 25455 20040 25467 20043
rect 25455 20012 26004 20040
rect 25455 20009 25467 20012
rect 25409 20003 25467 20009
rect 16224 19944 16804 19972
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15396 19876 15516 19904
rect 15580 19876 15945 19904
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19805 9643 19839
rect 9585 19799 9643 19805
rect 8389 19771 8447 19777
rect 8389 19737 8401 19771
rect 8435 19768 8447 19771
rect 9416 19768 9444 19799
rect 8435 19740 9444 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 8938 19700 8944 19712
rect 8312 19672 8944 19700
rect 7340 19660 7346 19672
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 9600 19700 9628 19799
rect 11330 19796 11336 19848
rect 11388 19796 11394 19848
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19836 14979 19839
rect 15378 19836 15384 19848
rect 14967 19808 15384 19836
rect 14967 19805 14979 19808
rect 14921 19799 14979 19805
rect 11793 19771 11851 19777
rect 11793 19737 11805 19771
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 9088 19672 9628 19700
rect 11241 19703 11299 19709
rect 9088 19660 9094 19672
rect 11241 19669 11253 19703
rect 11287 19700 11299 19703
rect 11808 19700 11836 19731
rect 12802 19728 12808 19780
rect 12860 19728 12866 19780
rect 14844 19768 14872 19799
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 15488 19845 15516 19876
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 15933 19867 15991 19873
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15562 19796 15568 19848
rect 15620 19796 15626 19848
rect 15746 19796 15752 19848
rect 15804 19796 15810 19848
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 16224 19836 16252 19944
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 18340 19904 18368 20000
rect 25976 19984 26004 20012
rect 18874 19932 18880 19984
rect 18932 19972 18938 19984
rect 19521 19975 19579 19981
rect 19521 19972 19533 19975
rect 18932 19944 19533 19972
rect 18932 19932 18938 19944
rect 19521 19941 19533 19944
rect 19567 19972 19579 19975
rect 20622 19972 20628 19984
rect 19567 19944 20628 19972
rect 19567 19941 19579 19944
rect 19521 19935 19579 19941
rect 20622 19932 20628 19944
rect 20680 19972 20686 19984
rect 20809 19975 20867 19981
rect 20809 19972 20821 19975
rect 20680 19944 20821 19972
rect 20680 19932 20686 19944
rect 20809 19941 20821 19944
rect 20855 19972 20867 19975
rect 21361 19975 21419 19981
rect 21361 19972 21373 19975
rect 20855 19944 21373 19972
rect 20855 19941 20867 19944
rect 20809 19935 20867 19941
rect 21361 19941 21373 19944
rect 21407 19941 21419 19975
rect 21361 19935 21419 19941
rect 25958 19932 25964 19984
rect 26016 19932 26022 19984
rect 18509 19907 18567 19913
rect 18509 19904 18521 19907
rect 16356 19876 16712 19904
rect 18340 19876 18521 19904
rect 16356 19864 16362 19876
rect 16172 19808 16252 19836
rect 16485 19839 16543 19845
rect 16172 19796 16178 19808
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 16531 19808 16620 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 16592 19780 16620 19808
rect 14844 19740 16246 19768
rect 11287 19672 11836 19700
rect 11287 19669 11299 19672
rect 11241 19663 11299 19669
rect 13354 19660 13360 19712
rect 13412 19700 13418 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 13412 19672 15301 19700
rect 13412 19660 13418 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 15289 19663 15347 19669
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 16022 19700 16028 19712
rect 15436 19672 16028 19700
rect 15436 19660 15442 19672
rect 16022 19660 16028 19672
rect 16080 19700 16086 19712
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 16080 19672 16129 19700
rect 16080 19660 16086 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16218 19700 16246 19740
rect 16574 19728 16580 19780
rect 16632 19728 16638 19780
rect 16684 19768 16712 19876
rect 18509 19873 18521 19876
rect 18555 19904 18567 19907
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 18555 19876 19257 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 19245 19873 19257 19876
rect 19291 19904 19303 19907
rect 19334 19904 19340 19916
rect 19291 19876 19340 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19904 21603 19907
rect 21591 19876 21864 19904
rect 21591 19873 21603 19876
rect 21545 19867 21603 19873
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 16777 19771 16835 19777
rect 16777 19768 16789 19771
rect 16684 19740 16789 19768
rect 16777 19737 16789 19740
rect 16823 19737 16835 19771
rect 19352 19768 19380 19864
rect 19720 19836 19748 19867
rect 21836 19845 21864 19876
rect 24118 19864 24124 19916
rect 24176 19904 24182 19916
rect 24670 19904 24676 19916
rect 24176 19876 24676 19904
rect 24176 19864 24182 19876
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19720 19808 19993 19836
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 19981 19799 20039 19805
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19836 24639 19839
rect 24854 19836 24860 19848
rect 24627 19808 24860 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 25225 19839 25283 19845
rect 25225 19805 25237 19839
rect 25271 19836 25283 19839
rect 26050 19836 26056 19848
rect 25271 19808 26056 19836
rect 25271 19805 25283 19808
rect 25225 19799 25283 19805
rect 26050 19796 26056 19808
rect 26108 19796 26114 19848
rect 20533 19771 20591 19777
rect 20533 19768 20545 19771
rect 19352 19740 20545 19768
rect 16777 19731 16835 19737
rect 20533 19737 20545 19740
rect 20579 19768 20591 19771
rect 21085 19771 21143 19777
rect 21085 19768 21097 19771
rect 20579 19740 21097 19768
rect 20579 19737 20591 19740
rect 20533 19731 20591 19737
rect 21085 19737 21097 19740
rect 21131 19737 21143 19771
rect 21085 19731 21143 19737
rect 23842 19728 23848 19780
rect 23900 19728 23906 19780
rect 23937 19771 23995 19777
rect 23937 19737 23949 19771
rect 23983 19768 23995 19771
rect 23983 19740 25268 19768
rect 23983 19737 23995 19740
rect 23937 19731 23995 19737
rect 25240 19712 25268 19740
rect 16945 19703 17003 19709
rect 16945 19700 16957 19703
rect 16218 19672 16957 19700
rect 16117 19663 16175 19669
rect 16945 19669 16957 19672
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 18046 19660 18052 19712
rect 18104 19660 18110 19712
rect 18969 19703 19027 19709
rect 18969 19669 18981 19703
rect 19015 19700 19027 19703
rect 19610 19700 19616 19712
rect 19015 19672 19616 19700
rect 19015 19669 19027 19672
rect 18969 19663 19027 19669
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 19794 19660 19800 19712
rect 19852 19660 19858 19712
rect 20990 19660 20996 19712
rect 21048 19660 21054 19712
rect 21542 19660 21548 19712
rect 21600 19700 21606 19712
rect 21637 19703 21695 19709
rect 21637 19700 21649 19703
rect 21600 19672 21649 19700
rect 21600 19660 21606 19672
rect 21637 19669 21649 19672
rect 21683 19669 21695 19703
rect 21637 19663 21695 19669
rect 23106 19660 23112 19712
rect 23164 19700 23170 19712
rect 23477 19703 23535 19709
rect 23477 19700 23489 19703
rect 23164 19672 23489 19700
rect 23164 19660 23170 19672
rect 23477 19669 23489 19672
rect 23523 19669 23535 19703
rect 23477 19663 23535 19669
rect 24394 19660 24400 19712
rect 24452 19660 24458 19712
rect 25222 19660 25228 19712
rect 25280 19660 25286 19712
rect 1104 19610 25852 19632
rect 1104 19558 4703 19610
rect 4755 19558 4767 19610
rect 4819 19558 4831 19610
rect 4883 19558 4895 19610
rect 4947 19558 4959 19610
rect 5011 19558 10890 19610
rect 10942 19558 10954 19610
rect 11006 19558 11018 19610
rect 11070 19558 11082 19610
rect 11134 19558 11146 19610
rect 11198 19558 17077 19610
rect 17129 19558 17141 19610
rect 17193 19558 17205 19610
rect 17257 19558 17269 19610
rect 17321 19558 17333 19610
rect 17385 19558 23264 19610
rect 23316 19558 23328 19610
rect 23380 19558 23392 19610
rect 23444 19558 23456 19610
rect 23508 19558 23520 19610
rect 23572 19558 25852 19610
rect 1104 19536 25852 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 2409 19499 2467 19505
rect 2409 19496 2421 19499
rect 2096 19468 2421 19496
rect 2096 19456 2102 19468
rect 2409 19465 2421 19468
rect 2455 19465 2467 19499
rect 2409 19459 2467 19465
rect 2590 19456 2596 19508
rect 2648 19456 2654 19508
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 2740 19468 4292 19496
rect 2740 19456 2746 19468
rect 1486 19320 1492 19372
rect 1544 19320 1550 19372
rect 1946 19320 1952 19372
rect 2004 19320 2010 19372
rect 2608 19369 2636 19456
rect 2700 19369 2728 19456
rect 3510 19388 3516 19440
rect 3568 19388 3574 19440
rect 4264 19428 4292 19468
rect 4338 19456 4344 19508
rect 4396 19496 4402 19508
rect 4396 19468 5028 19496
rect 4396 19456 4402 19468
rect 4430 19428 4436 19440
rect 4264 19400 4436 19428
rect 4430 19388 4436 19400
rect 4488 19388 4494 19440
rect 4522 19388 4528 19440
rect 4580 19428 4586 19440
rect 4580 19400 4844 19428
rect 4580 19388 4586 19400
rect 4816 19372 4844 19400
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19329 2651 19363
rect 2593 19323 2651 19329
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19329 2743 19363
rect 2685 19323 2743 19329
rect 4356 19332 4568 19360
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3602 19292 3608 19304
rect 3007 19264 3608 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3602 19252 3608 19264
rect 3660 19252 3666 19304
rect 1854 19184 1860 19236
rect 1912 19224 1918 19236
rect 1912 19196 2268 19224
rect 1912 19184 1918 19196
rect 2130 19116 2136 19168
rect 2188 19116 2194 19168
rect 2240 19156 2268 19196
rect 4356 19156 4384 19332
rect 4540 19304 4568 19332
rect 4798 19320 4804 19372
rect 4856 19320 4862 19372
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19261 4491 19295
rect 4433 19255 4491 19261
rect 4448 19224 4476 19255
rect 4522 19252 4528 19304
rect 4580 19252 4586 19304
rect 4614 19224 4620 19236
rect 4448 19196 4620 19224
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 5000 19224 5028 19468
rect 6454 19456 6460 19508
rect 6512 19456 6518 19508
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 7650 19496 7656 19508
rect 6963 19468 7656 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8352 19468 9413 19496
rect 8352 19456 8358 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10744 19468 10977 19496
rect 10744 19456 10750 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 12345 19499 12403 19505
rect 12345 19465 12357 19499
rect 12391 19496 12403 19499
rect 13078 19496 13084 19508
rect 12391 19468 13084 19496
rect 12391 19465 12403 19468
rect 12345 19459 12403 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13262 19456 13268 19508
rect 13320 19456 13326 19508
rect 14476 19468 17724 19496
rect 5902 19428 5908 19440
rect 5092 19400 5908 19428
rect 5092 19369 5120 19400
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5258 19320 5264 19372
rect 5316 19320 5322 19372
rect 5350 19320 5356 19372
rect 5408 19320 5414 19372
rect 6472 19369 6500 19456
rect 6549 19431 6607 19437
rect 6549 19397 6561 19431
rect 6595 19428 6607 19431
rect 6595 19400 6868 19428
rect 6595 19397 6607 19400
rect 6549 19391 6607 19397
rect 6840 19372 6868 19400
rect 7190 19388 7196 19440
rect 7248 19428 7254 19440
rect 7929 19431 7987 19437
rect 7929 19428 7941 19431
rect 7248 19400 7941 19428
rect 7248 19388 7254 19400
rect 7929 19397 7941 19400
rect 7975 19397 7987 19431
rect 7929 19391 7987 19397
rect 8570 19388 8576 19440
rect 8628 19388 8634 19440
rect 12710 19388 12716 19440
rect 12768 19388 12774 19440
rect 12805 19431 12863 19437
rect 12805 19397 12817 19431
rect 12851 19428 12863 19431
rect 14476 19428 14504 19468
rect 12851 19400 14504 19428
rect 14553 19431 14611 19437
rect 12851 19397 12863 19400
rect 12805 19391 12863 19397
rect 14553 19397 14565 19431
rect 14599 19428 14611 19431
rect 14826 19428 14832 19440
rect 14599 19400 14832 19428
rect 14599 19397 14611 19400
rect 14553 19391 14611 19397
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 15562 19388 15568 19440
rect 15620 19428 15626 19440
rect 15620 19400 16344 19428
rect 15620 19388 15626 19400
rect 5537 19363 5595 19369
rect 5537 19329 5549 19363
rect 5583 19360 5595 19363
rect 6457 19363 6515 19369
rect 5583 19332 6408 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 6380 19292 6408 19332
rect 6457 19329 6469 19363
rect 6503 19329 6515 19363
rect 6457 19323 6515 19329
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 6914 19320 6920 19372
rect 6972 19320 6978 19372
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7098 19360 7104 19372
rect 7055 19332 7104 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7098 19320 7104 19332
rect 7156 19360 7162 19372
rect 7156 19332 7512 19360
rect 7156 19320 7162 19332
rect 6932 19292 6960 19320
rect 6380 19264 6960 19292
rect 7484 19292 7512 19332
rect 7558 19320 7564 19372
rect 7616 19360 7622 19372
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 7616 19332 7665 19360
rect 7616 19320 7622 19332
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 10980 19332 11192 19360
rect 8386 19292 8392 19304
rect 7484 19264 8392 19292
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 9122 19292 9128 19304
rect 8536 19264 9128 19292
rect 8536 19252 8542 19264
rect 9122 19252 9128 19264
rect 9180 19292 9186 19304
rect 10980 19292 11008 19332
rect 9180 19264 11008 19292
rect 11057 19295 11115 19301
rect 9180 19252 9186 19264
rect 11057 19261 11069 19295
rect 11103 19261 11115 19295
rect 11164 19292 11192 19332
rect 12728 19358 12756 19388
rect 16316 19372 16344 19400
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 17034 19428 17040 19440
rect 16632 19400 17040 19428
rect 16632 19388 16638 19400
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 12820 19358 12940 19360
rect 12728 19332 12940 19358
rect 12728 19330 12848 19332
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 11164 19264 11253 19292
rect 11057 19255 11115 19261
rect 11241 19261 11253 19264
rect 11287 19292 11299 19295
rect 12342 19292 12348 19304
rect 11287 19264 12348 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 11072 19224 11100 19255
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 11606 19224 11612 19236
rect 5000 19196 5212 19224
rect 11072 19196 11612 19224
rect 5184 19168 5212 19196
rect 11606 19184 11612 19196
rect 11664 19224 11670 19236
rect 12452 19224 12480 19255
rect 12618 19252 12624 19304
rect 12676 19252 12682 19304
rect 12912 19301 12940 19332
rect 12986 19320 12992 19372
rect 13044 19358 13050 19372
rect 13081 19363 13139 19369
rect 13081 19358 13093 19363
rect 13044 19330 13093 19358
rect 13044 19320 13050 19330
rect 13081 19329 13093 19330
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 14240 19332 15301 19360
rect 14240 19320 14246 19332
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15436 19332 16037 19360
rect 15436 19320 15442 19332
rect 16025 19329 16037 19332
rect 16071 19329 16083 19363
rect 16025 19323 16083 19329
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 16172 19332 16221 19360
rect 16172 19320 16178 19332
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 16298 19320 16304 19372
rect 16356 19320 16362 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16776 19332 16865 19360
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 14366 19292 14372 19304
rect 12897 19255 12955 19261
rect 13004 19264 14372 19292
rect 12802 19224 12808 19236
rect 11664 19196 12388 19224
rect 12452 19196 12808 19224
rect 11664 19184 11670 19196
rect 2240 19128 4384 19156
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 4893 19159 4951 19165
rect 4893 19156 4905 19159
rect 4580 19128 4905 19156
rect 4580 19116 4586 19128
rect 4893 19125 4905 19128
rect 4939 19125 4951 19159
rect 4893 19119 4951 19125
rect 5166 19116 5172 19168
rect 5224 19116 5230 19168
rect 5810 19116 5816 19168
rect 5868 19116 5874 19168
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 9950 19156 9956 19168
rect 9824 19128 9956 19156
rect 9824 19116 9830 19128
rect 9950 19116 9956 19128
rect 10008 19116 10014 19168
rect 10597 19159 10655 19165
rect 10597 19125 10609 19159
rect 10643 19156 10655 19159
rect 10686 19156 10692 19168
rect 10643 19128 10692 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 11974 19116 11980 19168
rect 12032 19116 12038 19168
rect 12360 19156 12388 19196
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 13004 19156 13032 19264
rect 14366 19252 14372 19264
rect 14424 19292 14430 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14424 19264 14933 19292
rect 14424 19252 14430 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 15654 19292 15660 19304
rect 15252 19264 15660 19292
rect 15252 19252 15258 19264
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19292 15807 19295
rect 15930 19292 15936 19304
rect 15795 19264 15936 19292
rect 15795 19261 15807 19264
rect 15749 19255 15807 19261
rect 15930 19252 15936 19264
rect 15988 19292 15994 19304
rect 16776 19292 16804 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 15988 19264 16804 19292
rect 17696 19292 17724 19468
rect 17880 19468 19564 19496
rect 17880 19428 17908 19468
rect 17788 19400 17908 19428
rect 17788 19369 17816 19400
rect 18046 19388 18052 19440
rect 18104 19388 18110 19440
rect 19334 19428 19340 19440
rect 19274 19400 19340 19428
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 17773 19363 17831 19369
rect 17773 19329 17785 19363
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 18506 19292 18512 19304
rect 17696 19264 18512 19292
rect 15988 19252 15994 19264
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 19536 19292 19564 19468
rect 19794 19456 19800 19508
rect 19852 19456 19858 19508
rect 19886 19456 19892 19508
rect 19944 19496 19950 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 19944 19468 21373 19496
rect 19944 19456 19950 19468
rect 21361 19465 21373 19468
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 23106 19456 23112 19508
rect 23164 19456 23170 19508
rect 25222 19456 25228 19508
rect 25280 19496 25286 19508
rect 25280 19468 25820 19496
rect 25280 19456 25286 19468
rect 19812 19428 19840 19456
rect 19812 19400 20378 19428
rect 22186 19388 22192 19440
rect 22244 19388 22250 19440
rect 21634 19320 21640 19372
rect 21692 19320 21698 19372
rect 23124 19360 23152 19456
rect 23658 19388 23664 19440
rect 23716 19428 23722 19440
rect 23753 19431 23811 19437
rect 23753 19428 23765 19431
rect 23716 19400 23765 19428
rect 23716 19388 23722 19400
rect 23753 19397 23765 19400
rect 23799 19397 23811 19431
rect 23753 19391 23811 19397
rect 24394 19388 24400 19440
rect 24452 19388 24458 19440
rect 25792 19372 25820 19468
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23124 19332 23397 19360
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 23477 19363 23535 19369
rect 23477 19329 23489 19363
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19536 19264 19625 19292
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 14792 19196 15608 19224
rect 14792 19184 14798 19196
rect 12360 19128 13032 19156
rect 13078 19116 13084 19168
rect 13136 19116 13142 19168
rect 14918 19116 14924 19168
rect 14976 19156 14982 19168
rect 15197 19159 15255 19165
rect 15197 19156 15209 19159
rect 14976 19128 15209 19156
rect 14976 19116 14982 19128
rect 15197 19125 15209 19128
rect 15243 19125 15255 19159
rect 15197 19119 15255 19125
rect 15470 19116 15476 19168
rect 15528 19116 15534 19168
rect 15580 19156 15608 19196
rect 15838 19184 15844 19236
rect 15896 19184 15902 19236
rect 16666 19156 16672 19168
rect 15580 19128 16672 19156
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16758 19116 16764 19168
rect 16816 19116 16822 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 19484 19128 19533 19156
rect 19484 19116 19490 19128
rect 19521 19125 19533 19128
rect 19567 19125 19579 19159
rect 19628 19156 19656 19255
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 23014 19252 23020 19304
rect 23072 19292 23078 19304
rect 23492 19292 23520 19323
rect 25774 19320 25780 19372
rect 25832 19320 25838 19372
rect 23072 19264 23520 19292
rect 23072 19252 23078 19264
rect 21174 19184 21180 19236
rect 21232 19224 21238 19236
rect 21453 19227 21511 19233
rect 21453 19224 21465 19227
rect 21232 19196 21465 19224
rect 21232 19184 21238 19196
rect 21453 19193 21465 19196
rect 21499 19193 21511 19227
rect 21453 19187 21511 19193
rect 22373 19227 22431 19233
rect 22373 19193 22385 19227
rect 22419 19224 22431 19227
rect 23474 19224 23480 19236
rect 22419 19196 23480 19224
rect 22419 19193 22431 19196
rect 22373 19187 22431 19193
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 20530 19156 20536 19168
rect 19628 19128 20536 19156
rect 19521 19119 19579 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 23106 19116 23112 19168
rect 23164 19156 23170 19168
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 23164 19128 23213 19156
rect 23164 19116 23170 19128
rect 23201 19125 23213 19128
rect 23247 19125 23259 19159
rect 23201 19119 23259 19125
rect 1104 19066 25852 19088
rect 1104 19014 4043 19066
rect 4095 19014 4107 19066
rect 4159 19014 4171 19066
rect 4223 19014 4235 19066
rect 4287 19014 4299 19066
rect 4351 19014 10230 19066
rect 10282 19014 10294 19066
rect 10346 19014 10358 19066
rect 10410 19014 10422 19066
rect 10474 19014 10486 19066
rect 10538 19014 16417 19066
rect 16469 19014 16481 19066
rect 16533 19014 16545 19066
rect 16597 19014 16609 19066
rect 16661 19014 16673 19066
rect 16725 19014 22604 19066
rect 22656 19014 22668 19066
rect 22720 19014 22732 19066
rect 22784 19014 22796 19066
rect 22848 19014 22860 19066
rect 22912 19014 25852 19066
rect 1104 18992 25852 19014
rect 3786 18912 3792 18964
rect 3844 18912 3850 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 4890 18952 4896 18964
rect 4396 18924 4896 18952
rect 4396 18912 4402 18924
rect 4890 18912 4896 18924
rect 4948 18952 4954 18964
rect 5074 18952 5080 18964
rect 4948 18924 5080 18952
rect 4948 18912 4954 18924
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 5350 18912 5356 18964
rect 5408 18952 5414 18964
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 5408 18924 6469 18952
rect 5408 18912 5414 18924
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6457 18915 6515 18921
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 8018 18952 8024 18964
rect 6696 18924 8024 18952
rect 6696 18912 6702 18924
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 8128 18924 8493 18952
rect 4246 18884 4252 18896
rect 3620 18856 4252 18884
rect 3620 18828 3648 18856
rect 4246 18844 4252 18856
rect 4304 18884 4310 18896
rect 4304 18856 4844 18884
rect 4304 18844 4310 18856
rect 3602 18776 3608 18828
rect 3660 18776 3666 18828
rect 4338 18776 4344 18828
rect 4396 18776 4402 18828
rect 4816 18816 4844 18856
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 5629 18887 5687 18893
rect 5629 18884 5641 18887
rect 5316 18856 5641 18884
rect 5316 18844 5322 18856
rect 5629 18853 5641 18856
rect 5675 18853 5687 18887
rect 5629 18847 5687 18853
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 7374 18884 7380 18896
rect 5868 18856 7380 18884
rect 5868 18844 5874 18856
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 7650 18844 7656 18896
rect 7708 18884 7714 18896
rect 8128 18884 8156 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 9766 18952 9772 18964
rect 9548 18924 9772 18952
rect 9548 18912 9554 18924
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 11606 18912 11612 18964
rect 11664 18912 11670 18964
rect 14182 18912 14188 18964
rect 14240 18912 14246 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 14516 18924 14565 18952
rect 14516 18912 14522 18924
rect 14553 18921 14565 18924
rect 14599 18952 14611 18955
rect 14734 18952 14740 18964
rect 14599 18924 14740 18952
rect 14599 18921 14611 18924
rect 14553 18915 14611 18921
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 15381 18955 15439 18961
rect 15381 18952 15393 18955
rect 15344 18924 15393 18952
rect 15344 18912 15350 18924
rect 15381 18921 15393 18924
rect 15427 18921 15439 18955
rect 15381 18915 15439 18921
rect 15838 18912 15844 18964
rect 15896 18912 15902 18964
rect 15930 18912 15936 18964
rect 15988 18912 15994 18964
rect 16025 18955 16083 18961
rect 16025 18921 16037 18955
rect 16071 18921 16083 18955
rect 16025 18915 16083 18921
rect 7708 18856 8156 18884
rect 7708 18844 7714 18856
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 8662 18884 8668 18896
rect 8352 18856 8668 18884
rect 8352 18844 8358 18856
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 13924 18856 14970 18884
rect 4816 18788 4936 18816
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 4614 18748 4620 18760
rect 4295 18720 4620 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4908 18757 4936 18788
rect 5184 18788 5764 18816
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18717 4951 18751
rect 4893 18711 4951 18717
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18748 5135 18751
rect 5184 18748 5212 18788
rect 5736 18760 5764 18788
rect 7834 18776 7840 18828
rect 7892 18816 7898 18828
rect 8478 18816 8484 18828
rect 7892 18788 8484 18816
rect 7892 18776 7898 18788
rect 8478 18776 8484 18788
rect 8536 18816 8542 18828
rect 9030 18816 9036 18828
rect 8536 18788 9036 18816
rect 8536 18776 8542 18788
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9646 18788 9873 18816
rect 5123 18720 5212 18748
rect 5123 18717 5135 18720
rect 5077 18711 5135 18717
rect 5718 18708 5724 18760
rect 5776 18708 5782 18760
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 6086 18748 6092 18760
rect 5951 18720 6092 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7558 18748 7564 18760
rect 6972 18720 7564 18748
rect 6972 18708 6978 18720
rect 7558 18708 7564 18720
rect 7616 18748 7622 18760
rect 9646 18748 9674 18788
rect 9861 18785 9873 18788
rect 9907 18816 9919 18819
rect 11330 18816 11336 18828
rect 9907 18788 11336 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 13924 18760 13952 18856
rect 14942 18825 14970 18856
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15565 18887 15623 18893
rect 15565 18884 15577 18887
rect 15528 18856 15577 18884
rect 15528 18844 15534 18856
rect 15565 18853 15577 18856
rect 15611 18853 15623 18887
rect 15565 18847 15623 18853
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18785 14979 18819
rect 14921 18779 14979 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 15948 18816 15976 18912
rect 15896 18788 15976 18816
rect 15896 18776 15902 18788
rect 7616 18720 9674 18748
rect 7616 18708 7622 18720
rect 11974 18708 11980 18760
rect 12032 18708 12038 18760
rect 13906 18708 13912 18760
rect 13964 18708 13970 18760
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 4154 18640 4160 18692
rect 4212 18680 4218 18692
rect 5350 18680 5356 18692
rect 4212 18652 5356 18680
rect 4212 18640 4218 18652
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 8021 18683 8079 18689
rect 8021 18649 8033 18683
rect 8067 18680 8079 18683
rect 9030 18680 9036 18692
rect 8067 18652 9036 18680
rect 8067 18649 8079 18652
rect 8021 18643 8079 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 10134 18640 10140 18692
rect 10192 18640 10198 18692
rect 10594 18640 10600 18692
rect 10652 18640 10658 18692
rect 14108 18680 14136 18711
rect 14642 18708 14648 18760
rect 14700 18708 14706 18760
rect 14829 18751 14887 18757
rect 14829 18717 14841 18751
rect 14875 18717 14887 18751
rect 14829 18711 14887 18717
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18748 15071 18751
rect 15102 18748 15108 18760
rect 15059 18720 15108 18748
rect 15059 18717 15071 18720
rect 15013 18711 15071 18717
rect 14734 18680 14740 18692
rect 11716 18652 12020 18680
rect 14108 18652 14740 18680
rect 4614 18572 4620 18624
rect 4672 18612 4678 18624
rect 4801 18615 4859 18621
rect 4801 18612 4813 18615
rect 4672 18584 4813 18612
rect 4672 18572 4678 18584
rect 4801 18581 4813 18584
rect 4847 18581 4859 18615
rect 4801 18575 4859 18581
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 11716 18612 11744 18652
rect 11992 18624 12020 18652
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 4948 18584 11744 18612
rect 4948 18572 4954 18584
rect 11790 18572 11796 18624
rect 11848 18572 11854 18624
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 14844 18612 14872 18711
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15194 18708 15200 18760
rect 15252 18708 15258 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 15562 18748 15568 18760
rect 15519 18720 15568 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 15746 18708 15752 18760
rect 15804 18708 15810 18760
rect 16040 18748 16068 18915
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 16485 18955 16543 18961
rect 16485 18952 16497 18955
rect 16356 18924 16497 18952
rect 16356 18912 16362 18924
rect 16485 18921 16497 18924
rect 16531 18921 16543 18955
rect 16485 18915 16543 18921
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18230 18952 18236 18964
rect 18187 18924 18236 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19392 18924 19533 18952
rect 19392 18912 19398 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 19886 18912 19892 18964
rect 19944 18912 19950 18964
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 24486 18952 24492 18964
rect 20036 18924 24492 18952
rect 20036 18912 20042 18924
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 24854 18912 24860 18964
rect 24912 18912 24918 18964
rect 25406 18912 25412 18964
rect 25464 18912 25470 18964
rect 17773 18887 17831 18893
rect 17773 18853 17785 18887
rect 17819 18884 17831 18887
rect 19245 18887 19303 18893
rect 17819 18856 18920 18884
rect 17819 18853 17831 18856
rect 17773 18847 17831 18853
rect 16209 18819 16267 18825
rect 16209 18785 16221 18819
rect 16255 18816 16267 18819
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 16255 18788 16804 18816
rect 16255 18785 16267 18788
rect 16209 18779 16267 18785
rect 16776 18760 16804 18788
rect 16960 18788 17877 18816
rect 15856 18720 16068 18748
rect 16301 18751 16359 18757
rect 14918 18640 14924 18692
rect 14976 18640 14982 18692
rect 15378 18640 15384 18692
rect 15436 18680 15442 18692
rect 15856 18680 15884 18720
rect 16301 18717 16313 18751
rect 16347 18748 16359 18751
rect 16482 18748 16488 18760
rect 16347 18720 16488 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16666 18748 16672 18760
rect 16623 18720 16672 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 16960 18757 16988 18788
rect 17865 18785 17877 18788
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17494 18748 17500 18760
rect 17175 18720 17500 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 18506 18708 18512 18760
rect 18564 18708 18570 18760
rect 18616 18757 18644 18856
rect 18782 18776 18788 18828
rect 18840 18776 18846 18828
rect 18892 18816 18920 18856
rect 19245 18853 19257 18887
rect 19291 18884 19303 18887
rect 19904 18884 19932 18912
rect 19291 18856 19932 18884
rect 19291 18853 19303 18856
rect 19245 18847 19303 18853
rect 23934 18844 23940 18896
rect 23992 18884 23998 18896
rect 24673 18887 24731 18893
rect 24673 18884 24685 18887
rect 23992 18856 24685 18884
rect 23992 18844 23998 18856
rect 24673 18853 24685 18856
rect 24719 18853 24731 18887
rect 24673 18847 24731 18853
rect 19334 18816 19340 18828
rect 18892 18788 19340 18816
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19610 18776 19616 18828
rect 19668 18776 19674 18828
rect 20530 18776 20536 18828
rect 20588 18816 20594 18828
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 20588 18788 20637 18816
rect 20588 18776 20594 18788
rect 20625 18785 20637 18788
rect 20671 18816 20683 18819
rect 20671 18788 23060 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18800 18748 18828 18776
rect 18800 18720 19334 18748
rect 18601 18711 18659 18717
rect 15436 18652 15884 18680
rect 16025 18683 16083 18689
rect 15436 18640 15442 18652
rect 16025 18649 16037 18683
rect 16071 18680 16083 18683
rect 16071 18652 16804 18680
rect 16071 18649 16083 18652
rect 16025 18643 16083 18649
rect 14936 18612 14964 18640
rect 14844 18584 14964 18612
rect 15102 18572 15108 18624
rect 15160 18612 15166 18624
rect 16669 18615 16727 18621
rect 16669 18612 16681 18615
rect 15160 18584 16681 18612
rect 15160 18572 15166 18584
rect 16669 18581 16681 18584
rect 16715 18581 16727 18615
rect 16776 18612 16804 18652
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17405 18683 17463 18689
rect 17405 18680 17417 18683
rect 16908 18652 17417 18680
rect 16908 18640 16914 18652
rect 17405 18649 17417 18652
rect 17451 18680 17463 18683
rect 17770 18680 17776 18692
rect 17451 18652 17776 18680
rect 17451 18649 17463 18652
rect 17405 18643 17463 18649
rect 17770 18640 17776 18652
rect 17828 18640 17834 18692
rect 19306 18680 19334 18720
rect 19426 18708 19432 18760
rect 19484 18708 19490 18760
rect 19628 18748 19656 18776
rect 23032 18760 23060 18788
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 23658 18816 23664 18828
rect 23532 18788 23664 18816
rect 23532 18776 23538 18788
rect 23658 18776 23664 18788
rect 23716 18816 23722 18828
rect 24397 18819 24455 18825
rect 24397 18816 24409 18819
rect 23716 18788 24409 18816
rect 23716 18776 23722 18788
rect 24397 18785 24409 18788
rect 24443 18785 24455 18819
rect 24397 18779 24455 18785
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19628 18720 19717 18748
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 23014 18708 23020 18760
rect 23072 18708 23078 18760
rect 25130 18708 25136 18760
rect 25188 18708 25194 18760
rect 25222 18708 25228 18760
rect 25280 18708 25286 18760
rect 19886 18680 19892 18692
rect 19306 18652 19892 18680
rect 19886 18640 19892 18652
rect 19944 18640 19950 18692
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 21174 18680 21180 18692
rect 20947 18652 21180 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 21542 18640 21548 18692
rect 21600 18640 21606 18692
rect 17034 18612 17040 18624
rect 16776 18584 17040 18612
rect 16669 18575 16727 18581
rect 17034 18572 17040 18584
rect 17092 18612 17098 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 17092 18584 17325 18612
rect 17092 18572 17098 18584
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 22278 18612 22284 18624
rect 17644 18584 22284 18612
rect 17644 18572 17650 18584
rect 22278 18572 22284 18584
rect 22336 18612 22342 18624
rect 22373 18615 22431 18621
rect 22373 18612 22385 18615
rect 22336 18584 22385 18612
rect 22336 18572 22342 18584
rect 22373 18581 22385 18584
rect 22419 18581 22431 18615
rect 22373 18575 22431 18581
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 1104 18522 25852 18544
rect 1104 18470 4703 18522
rect 4755 18470 4767 18522
rect 4819 18470 4831 18522
rect 4883 18470 4895 18522
rect 4947 18470 4959 18522
rect 5011 18470 10890 18522
rect 10942 18470 10954 18522
rect 11006 18470 11018 18522
rect 11070 18470 11082 18522
rect 11134 18470 11146 18522
rect 11198 18470 17077 18522
rect 17129 18470 17141 18522
rect 17193 18470 17205 18522
rect 17257 18470 17269 18522
rect 17321 18470 17333 18522
rect 17385 18470 23264 18522
rect 23316 18470 23328 18522
rect 23380 18470 23392 18522
rect 23444 18470 23456 18522
rect 23508 18470 23520 18522
rect 23572 18470 25852 18522
rect 1104 18448 25852 18470
rect 4522 18368 4528 18420
rect 4580 18408 4586 18420
rect 4580 18380 4660 18408
rect 4580 18368 4586 18380
rect 4632 18349 4660 18380
rect 7116 18380 7880 18408
rect 4617 18343 4675 18349
rect 4617 18309 4629 18343
rect 4663 18309 4675 18343
rect 6362 18340 6368 18352
rect 5842 18312 6368 18340
rect 4617 18303 4675 18309
rect 6362 18300 6368 18312
rect 6420 18300 6426 18352
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 3050 18272 3056 18284
rect 2363 18244 3056 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 7006 18232 7012 18284
rect 7064 18232 7070 18284
rect 4338 18164 4344 18216
rect 4396 18164 4402 18216
rect 7116 18204 7144 18380
rect 7285 18343 7343 18349
rect 7285 18309 7297 18343
rect 7331 18340 7343 18343
rect 7331 18312 7420 18340
rect 7331 18309 7343 18312
rect 7285 18303 7343 18309
rect 7190 18204 7196 18216
rect 4448 18176 7196 18204
rect 2222 18096 2228 18148
rect 2280 18136 2286 18148
rect 4448 18136 4476 18176
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7392 18204 7420 18312
rect 7852 18296 7880 18380
rect 8938 18368 8944 18420
rect 8996 18368 9002 18420
rect 9214 18368 9220 18420
rect 9272 18368 9278 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 10192 18380 10333 18408
rect 10192 18368 10198 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 10321 18371 10379 18377
rect 10686 18368 10692 18420
rect 10744 18368 10750 18420
rect 12802 18368 12808 18420
rect 12860 18408 12866 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 12860 18380 13277 18408
rect 12860 18368 12866 18380
rect 13265 18377 13277 18380
rect 13311 18408 13323 18411
rect 13906 18408 13912 18420
rect 13311 18380 13912 18408
rect 13311 18377 13323 18380
rect 13265 18371 13323 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14093 18411 14151 18417
rect 14093 18377 14105 18411
rect 14139 18408 14151 18411
rect 15746 18408 15752 18420
rect 14139 18380 15752 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 16482 18408 16488 18420
rect 15988 18380 16488 18408
rect 15988 18368 15994 18380
rect 16482 18368 16488 18380
rect 16540 18368 16546 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 19978 18408 19984 18420
rect 16724 18380 19984 18408
rect 16724 18368 16730 18380
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20990 18368 20996 18420
rect 21048 18368 21054 18420
rect 21634 18368 21640 18420
rect 21692 18408 21698 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 21692 18380 21833 18408
rect 21692 18368 21698 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 21821 18371 21879 18377
rect 22278 18368 22284 18420
rect 22336 18368 22342 18420
rect 23106 18368 23112 18420
rect 23164 18408 23170 18420
rect 23164 18380 23428 18408
rect 23164 18368 23170 18380
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18262 7527 18275
rect 7558 18262 7564 18284
rect 7515 18241 7564 18262
rect 7469 18235 7564 18241
rect 7484 18234 7564 18235
rect 7558 18232 7564 18234
rect 7616 18232 7622 18284
rect 7650 18232 7656 18284
rect 7708 18232 7714 18284
rect 7760 18281 7880 18296
rect 7745 18275 7880 18281
rect 7745 18241 7757 18275
rect 7791 18268 7880 18275
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 7791 18241 7803 18268
rect 7745 18235 7803 18241
rect 7944 18244 8585 18272
rect 7944 18204 7972 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 9232 18272 9260 18368
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9232 18244 10149 18272
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 10704 18272 10732 18368
rect 12434 18300 12440 18352
rect 12492 18300 12498 18352
rect 14642 18340 14648 18352
rect 14016 18312 14648 18340
rect 14016 18281 14044 18312
rect 14642 18300 14648 18312
rect 14700 18340 14706 18352
rect 15378 18340 15384 18352
rect 14700 18312 15384 18340
rect 14700 18300 14706 18312
rect 15378 18300 15384 18312
rect 15436 18300 15442 18352
rect 15470 18300 15476 18352
rect 15528 18300 15534 18352
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 16301 18343 16359 18349
rect 16301 18340 16313 18343
rect 15896 18312 16313 18340
rect 15896 18300 15902 18312
rect 16301 18309 16313 18312
rect 16347 18309 16359 18343
rect 16301 18303 16359 18309
rect 16390 18300 16396 18352
rect 16448 18340 16454 18352
rect 17402 18340 17408 18352
rect 16448 18312 17408 18340
rect 16448 18300 16454 18312
rect 17402 18300 17408 18312
rect 17460 18340 17466 18352
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 17460 18312 18245 18340
rect 17460 18300 17466 18312
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 10551 18244 10732 18272
rect 14001 18275 14059 18281
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 14001 18241 14013 18275
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 7392 18176 7972 18204
rect 7285 18167 7343 18173
rect 2280 18108 4476 18136
rect 2280 18096 2286 18108
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 2096 18040 2145 18068
rect 2096 18028 2102 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2133 18031 2191 18037
rect 6086 18028 6092 18080
rect 6144 18028 6150 18080
rect 7098 18028 7104 18080
rect 7156 18028 7162 18080
rect 7300 18068 7328 18167
rect 8018 18164 8024 18216
rect 8076 18164 8082 18216
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18173 8539 18207
rect 8680 18204 8708 18232
rect 9490 18204 9496 18216
rect 8680 18176 9496 18204
rect 8481 18167 8539 18173
rect 7469 18139 7527 18145
rect 7469 18105 7481 18139
rect 7515 18136 7527 18139
rect 8496 18136 8524 18167
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11388 18176 11529 18204
rect 11388 18164 11394 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 11790 18164 11796 18216
rect 11848 18164 11854 18216
rect 7515 18108 8524 18136
rect 14200 18136 14228 18235
rect 14366 18232 14372 18284
rect 14424 18232 14430 18284
rect 15102 18272 15108 18284
rect 15042 18244 15108 18272
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 14384 18204 14412 18232
rect 15212 18204 15240 18232
rect 14384 18176 15240 18204
rect 15488 18204 15516 18300
rect 15562 18232 15568 18284
rect 15620 18232 15626 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15764 18204 15792 18235
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16080 18244 16681 18272
rect 16080 18232 16086 18244
rect 16669 18241 16681 18244
rect 16715 18272 16727 18275
rect 17034 18272 17040 18284
rect 16715 18244 17040 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 17494 18272 17500 18284
rect 17175 18244 17500 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18272 17739 18275
rect 17770 18272 17776 18284
rect 17727 18244 17776 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 19334 18272 19340 18284
rect 17911 18244 19340 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20530 18272 20536 18284
rect 20027 18244 20536 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 21008 18272 21036 18368
rect 22189 18343 22247 18349
rect 22189 18309 22201 18343
rect 22235 18340 22247 18343
rect 23290 18340 23296 18352
rect 22235 18312 23296 18340
rect 22235 18309 22247 18312
rect 22189 18303 22247 18309
rect 23290 18300 23296 18312
rect 23348 18300 23354 18352
rect 23400 18349 23428 18380
rect 23385 18343 23443 18349
rect 23385 18309 23397 18343
rect 23431 18309 23443 18343
rect 24946 18340 24952 18352
rect 24610 18312 24952 18340
rect 23385 18303 23443 18309
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 25958 18340 25964 18352
rect 25516 18312 25964 18340
rect 25516 18281 25544 18312
rect 25958 18300 25964 18312
rect 26016 18300 26022 18352
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 21008 18244 21465 18272
rect 21453 18241 21465 18244
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 15488 18176 15792 18204
rect 14200 18108 15424 18136
rect 7515 18105 7527 18108
rect 7469 18099 7527 18105
rect 15396 18080 15424 18108
rect 7926 18068 7932 18080
rect 7300 18040 7932 18068
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 8110 18028 8116 18080
rect 8168 18028 8174 18080
rect 8294 18028 8300 18080
rect 8352 18028 8358 18080
rect 15378 18028 15384 18080
rect 15436 18028 15442 18080
rect 15764 18068 15792 18176
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 16816 18176 17417 18204
rect 16816 18164 16822 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 17512 18204 17540 18232
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17512 18176 18061 18204
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 15933 18139 15991 18145
rect 15933 18136 15945 18139
rect 15896 18108 15945 18136
rect 15896 18096 15902 18108
rect 15933 18105 15945 18108
rect 15979 18105 15991 18139
rect 17512 18136 17540 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18156 18176 22232 18204
rect 15933 18099 15991 18105
rect 16684 18108 17540 18136
rect 16684 18077 16712 18108
rect 17770 18096 17776 18148
rect 17828 18136 17834 18148
rect 18156 18136 18184 18176
rect 21634 18136 21640 18148
rect 17828 18108 18184 18136
rect 18524 18108 21640 18136
rect 17828 18096 17834 18108
rect 18524 18080 18552 18108
rect 21634 18096 21640 18108
rect 21692 18096 21698 18148
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 15764 18040 16681 18068
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17034 18028 17040 18080
rect 17092 18028 17098 18080
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 17221 18071 17279 18077
rect 17221 18068 17233 18071
rect 17184 18040 17233 18068
rect 17184 18028 17190 18040
rect 17221 18037 17233 18040
rect 17267 18037 17279 18071
rect 17221 18031 17279 18037
rect 17310 18028 17316 18080
rect 17368 18028 17374 18080
rect 18506 18028 18512 18080
rect 18564 18028 18570 18080
rect 21266 18028 21272 18080
rect 21324 18028 21330 18080
rect 22204 18068 22232 18176
rect 22370 18164 22376 18216
rect 22428 18164 22434 18216
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 23072 18176 23121 18204
rect 23072 18164 23078 18176
rect 23109 18173 23121 18176
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 24486 18068 24492 18080
rect 22204 18040 24492 18068
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 24854 18028 24860 18080
rect 24912 18028 24918 18080
rect 25314 18028 25320 18080
rect 25372 18028 25378 18080
rect 1104 17978 25852 18000
rect 1104 17926 4043 17978
rect 4095 17926 4107 17978
rect 4159 17926 4171 17978
rect 4223 17926 4235 17978
rect 4287 17926 4299 17978
rect 4351 17926 10230 17978
rect 10282 17926 10294 17978
rect 10346 17926 10358 17978
rect 10410 17926 10422 17978
rect 10474 17926 10486 17978
rect 10538 17926 16417 17978
rect 16469 17926 16481 17978
rect 16533 17926 16545 17978
rect 16597 17926 16609 17978
rect 16661 17926 16673 17978
rect 16725 17926 22604 17978
rect 22656 17926 22668 17978
rect 22720 17926 22732 17978
rect 22784 17926 22796 17978
rect 22848 17926 22860 17978
rect 22912 17926 25852 17978
rect 1104 17904 25852 17926
rect 4430 17824 4436 17876
rect 4488 17864 4494 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 4488 17836 6745 17864
rect 4488 17824 4494 17836
rect 6733 17833 6745 17836
rect 6779 17864 6791 17867
rect 6914 17864 6920 17876
rect 6779 17836 6920 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7558 17864 7564 17876
rect 7432 17836 7564 17864
rect 7432 17824 7438 17836
rect 7558 17824 7564 17836
rect 7616 17864 7622 17876
rect 8110 17864 8116 17876
rect 7616 17836 8116 17864
rect 7616 17824 7622 17836
rect 8110 17824 8116 17836
rect 8168 17864 8174 17876
rect 8168 17836 8800 17864
rect 8168 17824 8174 17836
rect 8665 17799 8723 17805
rect 8665 17796 8677 17799
rect 7668 17768 8677 17796
rect 1670 17688 1676 17740
rect 1728 17688 1734 17740
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2038 17728 2044 17740
rect 1995 17700 2044 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 3421 17731 3479 17737
rect 3421 17697 3433 17731
rect 3467 17728 3479 17731
rect 3694 17728 3700 17740
rect 3467 17700 3700 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 3694 17688 3700 17700
rect 3752 17728 3758 17740
rect 4249 17731 4307 17737
rect 4249 17728 4261 17731
rect 3752 17700 4016 17728
rect 3752 17688 3758 17700
rect 3988 17669 4016 17700
rect 4080 17700 4261 17728
rect 4080 17672 4108 17700
rect 4249 17697 4261 17700
rect 4295 17697 4307 17731
rect 7668 17728 7696 17768
rect 8665 17765 8677 17768
rect 8711 17765 8723 17799
rect 8772 17796 8800 17836
rect 9030 17824 9036 17876
rect 9088 17824 9094 17876
rect 9953 17867 10011 17873
rect 9953 17864 9965 17867
rect 9140 17836 9965 17864
rect 9140 17796 9168 17836
rect 9953 17833 9965 17836
rect 9999 17833 10011 17867
rect 9953 17827 10011 17833
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 13262 17864 13268 17876
rect 12023 17836 13268 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13906 17824 13912 17876
rect 13964 17824 13970 17876
rect 15562 17824 15568 17876
rect 15620 17864 15626 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 15620 17836 15669 17864
rect 15620 17824 15626 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 15930 17864 15936 17876
rect 15657 17827 15715 17833
rect 15764 17836 15936 17864
rect 9769 17799 9827 17805
rect 9769 17796 9781 17799
rect 8772 17768 9168 17796
rect 9508 17768 9781 17796
rect 8665 17759 8723 17765
rect 4249 17691 4307 17697
rect 7024 17700 7696 17728
rect 7024 17672 7052 17700
rect 7668 17672 7696 17700
rect 7926 17688 7932 17740
rect 7984 17728 7990 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 7984 17700 8432 17728
rect 7984 17688 7990 17700
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 4062 17620 4068 17672
rect 4120 17620 4126 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 4172 17592 4200 17623
rect 5258 17620 5264 17672
rect 5316 17620 5322 17672
rect 7006 17620 7012 17672
rect 7064 17620 7070 17672
rect 7374 17620 7380 17672
rect 7432 17620 7438 17672
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8294 17660 8300 17672
rect 8159 17632 8300 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 2280 17564 2438 17592
rect 3988 17564 4200 17592
rect 2280 17552 2286 17564
rect 3988 17536 4016 17564
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 2924 17496 3801 17524
rect 2924 17484 2930 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 3789 17487 3847 17493
rect 3970 17484 3976 17536
rect 4028 17484 4034 17536
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7852 17524 7880 17623
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 8404 17592 8432 17700
rect 8496 17700 9413 17728
rect 8496 17669 8524 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 8570 17620 8576 17672
rect 8628 17620 8634 17672
rect 8754 17662 8760 17672
rect 8680 17634 8760 17662
rect 8680 17592 8708 17634
rect 8754 17620 8760 17634
rect 8812 17620 8818 17672
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 8404 17564 8708 17592
rect 8956 17592 8984 17623
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9508 17660 9536 17768
rect 9769 17765 9781 17768
rect 9815 17765 9827 17799
rect 9769 17759 9827 17765
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 9732 17700 11805 17728
rect 9732 17688 9738 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 13924 17728 13952 17824
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 13924 17700 14657 17728
rect 11793 17691 11851 17697
rect 14645 17697 14657 17700
rect 14691 17728 14703 17731
rect 14734 17728 14740 17740
rect 14691 17700 14740 17728
rect 14691 17697 14703 17700
rect 14645 17691 14703 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 14826 17688 14832 17740
rect 14884 17728 14890 17740
rect 15470 17728 15476 17740
rect 14884 17700 15476 17728
rect 14884 17688 14890 17700
rect 9088 17632 9720 17660
rect 9088 17620 9094 17632
rect 9692 17604 9720 17632
rect 10778 17620 10784 17672
rect 10836 17620 10842 17672
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12023 17632 14412 17660
rect 15120 17646 15148 17700
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 9490 17592 9496 17604
rect 8956 17564 9496 17592
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 9674 17552 9680 17604
rect 9732 17552 9738 17604
rect 11698 17552 11704 17604
rect 11756 17552 11762 17604
rect 7926 17524 7932 17536
rect 7156 17496 7932 17524
rect 7156 17484 7162 17496
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8444 17496 8493 17524
rect 8444 17484 8450 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 8481 17487 8539 17493
rect 12161 17527 12219 17533
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 13722 17524 13728 17536
rect 12207 17496 13728 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 14384 17524 14412 17632
rect 15304 17632 15577 17660
rect 14458 17552 14464 17604
rect 14516 17592 14522 17604
rect 15304 17592 15332 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 14516 17564 15332 17592
rect 14516 17552 14522 17564
rect 15378 17552 15384 17604
rect 15436 17592 15442 17604
rect 15473 17595 15531 17601
rect 15473 17592 15485 17595
rect 15436 17564 15485 17592
rect 15436 17552 15442 17564
rect 15473 17561 15485 17564
rect 15519 17592 15531 17595
rect 15764 17592 15792 17836
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 19245 17867 19303 17873
rect 19245 17833 19257 17867
rect 19291 17864 19303 17867
rect 19426 17864 19432 17876
rect 19291 17836 19432 17864
rect 19291 17833 19303 17836
rect 19245 17827 19303 17833
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 19668 17836 22094 17864
rect 19668 17824 19674 17836
rect 17310 17796 17316 17808
rect 15948 17768 17316 17796
rect 15948 17669 15976 17768
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 22066 17796 22094 17836
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 23109 17867 23167 17873
rect 23109 17864 23121 17867
rect 22520 17836 23121 17864
rect 22520 17824 22526 17836
rect 23109 17833 23121 17836
rect 23155 17833 23167 17867
rect 23109 17827 23167 17833
rect 23198 17824 23204 17876
rect 23256 17824 23262 17876
rect 24121 17867 24179 17873
rect 24121 17833 24133 17867
rect 24167 17864 24179 17867
rect 25130 17864 25136 17876
rect 24167 17836 25136 17864
rect 24167 17833 24179 17836
rect 24121 17827 24179 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 23216 17796 23244 17824
rect 23569 17799 23627 17805
rect 23569 17796 23581 17799
rect 22066 17768 23152 17796
rect 23216 17768 23581 17796
rect 16025 17731 16083 17737
rect 16025 17697 16037 17731
rect 16071 17728 16083 17731
rect 16071 17700 16344 17728
rect 16071 17697 16083 17700
rect 16025 17691 16083 17697
rect 16316 17672 16344 17700
rect 19886 17688 19892 17740
rect 19944 17728 19950 17740
rect 22186 17728 22192 17740
rect 19944 17700 22192 17728
rect 19944 17688 19950 17700
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 15519 17564 15792 17592
rect 15856 17592 15884 17623
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 17034 17620 17040 17672
rect 17092 17620 17098 17672
rect 20530 17620 20536 17672
rect 20588 17620 20594 17672
rect 23124 17669 23152 17768
rect 23569 17765 23581 17768
rect 23615 17765 23627 17799
rect 23569 17759 23627 17765
rect 23934 17756 23940 17808
rect 23992 17756 23998 17808
rect 24394 17756 24400 17808
rect 24452 17756 24458 17808
rect 24670 17756 24676 17808
rect 24728 17796 24734 17808
rect 24728 17768 24992 17796
rect 24728 17756 24734 17768
rect 23201 17731 23259 17737
rect 23201 17697 23213 17731
rect 23247 17697 23259 17731
rect 23201 17691 23259 17697
rect 22373 17663 22431 17669
rect 22373 17660 22385 17663
rect 22296 17632 22385 17660
rect 17052 17592 17080 17620
rect 15856 17564 17080 17592
rect 19705 17595 19763 17601
rect 15519 17561 15531 17564
rect 15473 17555 15531 17561
rect 19705 17561 19717 17595
rect 19751 17592 19763 17595
rect 19794 17592 19800 17604
rect 19751 17564 19800 17592
rect 19751 17561 19763 17564
rect 19705 17555 19763 17561
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 20806 17552 20812 17604
rect 20864 17552 20870 17604
rect 21266 17552 21272 17604
rect 21324 17552 21330 17604
rect 16022 17524 16028 17536
rect 14384 17496 16028 17524
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 16114 17484 16120 17536
rect 16172 17484 16178 17536
rect 19610 17484 19616 17536
rect 19668 17484 19674 17536
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 22296 17533 22324 17632
rect 22373 17629 22385 17632
rect 22419 17629 22431 17663
rect 22373 17623 22431 17629
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 22830 17552 22836 17604
rect 22888 17592 22894 17604
rect 23216 17592 23244 17691
rect 23658 17688 23664 17740
rect 23716 17688 23722 17740
rect 24118 17688 24124 17740
rect 24176 17728 24182 17740
rect 24854 17728 24860 17740
rect 24176 17700 24860 17728
rect 24176 17688 24182 17700
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 24964 17737 24992 17768
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 23348 17632 23397 17660
rect 23348 17620 23354 17632
rect 23385 17629 23397 17632
rect 23431 17660 23443 17663
rect 23431 17632 23796 17660
rect 23431 17629 23443 17632
rect 23385 17623 23443 17629
rect 23768 17592 23796 17632
rect 24026 17620 24032 17672
rect 24084 17660 24090 17672
rect 24765 17663 24823 17669
rect 24765 17660 24777 17663
rect 24084 17632 24777 17660
rect 24084 17620 24090 17632
rect 24765 17629 24777 17632
rect 24811 17629 24823 17663
rect 24765 17623 24823 17629
rect 22888 17564 23704 17592
rect 23768 17564 25912 17592
rect 22888 17552 22894 17564
rect 22281 17527 22339 17533
rect 22281 17524 22293 17527
rect 21876 17496 22293 17524
rect 21876 17484 21882 17496
rect 22281 17493 22293 17496
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22704 17496 23029 17524
rect 22704 17484 22710 17496
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 23676 17524 23704 17564
rect 25130 17524 25136 17536
rect 23676 17496 25136 17524
rect 23017 17487 23075 17493
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 1104 17434 25852 17456
rect 1104 17382 4703 17434
rect 4755 17382 4767 17434
rect 4819 17382 4831 17434
rect 4883 17382 4895 17434
rect 4947 17382 4959 17434
rect 5011 17382 10890 17434
rect 10942 17382 10954 17434
rect 11006 17382 11018 17434
rect 11070 17382 11082 17434
rect 11134 17382 11146 17434
rect 11198 17382 17077 17434
rect 17129 17382 17141 17434
rect 17193 17382 17205 17434
rect 17257 17382 17269 17434
rect 17321 17382 17333 17434
rect 17385 17382 23264 17434
rect 23316 17382 23328 17434
rect 23380 17382 23392 17434
rect 23444 17382 23456 17434
rect 23508 17382 23520 17434
rect 23572 17382 25852 17434
rect 1104 17360 25852 17382
rect 2222 17280 2228 17332
rect 2280 17280 2286 17332
rect 2866 17280 2872 17332
rect 2924 17280 2930 17332
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 3694 17280 3700 17332
rect 3752 17280 3758 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3804 17292 4077 17320
rect 1394 17144 1400 17196
rect 1452 17144 1458 17196
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2774 17184 2780 17196
rect 2547 17156 2780 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1688 17116 1716 17147
rect 992 17088 1716 17116
rect 992 17076 998 17088
rect 1578 17008 1584 17060
rect 1636 17008 1642 17060
rect 2424 17048 2452 17147
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 2884 17193 2912 17280
rect 3712 17193 3740 17280
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 3697 17187 3755 17193
rect 2869 17147 2927 17153
rect 3068 17156 3648 17184
rect 2792 17116 2820 17144
rect 3068 17116 3096 17156
rect 2792 17088 3096 17116
rect 3142 17076 3148 17128
rect 3200 17076 3206 17128
rect 3620 17116 3648 17156
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3804 17116 3832 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 4065 17283 4123 17289
rect 4430 17280 4436 17332
rect 4488 17280 4494 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 5960 17292 6653 17320
rect 5960 17280 5966 17292
rect 6641 17289 6653 17292
rect 6687 17289 6699 17323
rect 6641 17283 6699 17289
rect 7377 17323 7435 17329
rect 7377 17289 7389 17323
rect 7423 17320 7435 17323
rect 8570 17320 8576 17332
rect 7423 17292 8576 17320
rect 7423 17289 7435 17292
rect 7377 17283 7435 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 8754 17280 8760 17332
rect 8812 17320 8818 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 8812 17292 9137 17320
rect 8812 17280 8818 17292
rect 9125 17289 9137 17292
rect 9171 17289 9183 17323
rect 9125 17283 9183 17289
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 12434 17320 12440 17332
rect 10919 17292 12440 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15654 17320 15660 17332
rect 14792 17292 15660 17320
rect 14792 17280 14798 17292
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16264 17292 16957 17320
rect 16264 17280 16270 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 16945 17283 17003 17289
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20864 17292 21097 17320
rect 20864 17280 20870 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 21085 17283 21143 17289
rect 22281 17323 22339 17329
rect 22281 17289 22293 17323
rect 22327 17320 22339 17323
rect 22646 17320 22652 17332
rect 22327 17292 22652 17320
rect 22327 17289 22339 17292
rect 22281 17283 22339 17289
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 22830 17280 22836 17332
rect 22888 17280 22894 17332
rect 23106 17280 23112 17332
rect 23164 17280 23170 17332
rect 24394 17320 24400 17332
rect 23584 17292 24400 17320
rect 4448 17252 4476 17280
rect 4356 17224 4476 17252
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 4062 17184 4068 17196
rect 3927 17156 4068 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4356 17193 4384 17224
rect 4614 17212 4620 17264
rect 4672 17212 4678 17264
rect 5994 17252 6000 17264
rect 5842 17224 6000 17252
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 7190 17212 7196 17264
rect 7248 17252 7254 17264
rect 7248 17224 8248 17252
rect 7248 17212 7254 17224
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 6963 17156 7604 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 3620 17088 3832 17116
rect 4080 17116 4108 17144
rect 6089 17119 6147 17125
rect 6089 17116 6101 17119
rect 4080 17088 6101 17116
rect 3712 17060 3740 17088
rect 5736 17060 5764 17088
rect 6089 17085 6101 17088
rect 6135 17116 6147 17119
rect 6380 17116 6408 17147
rect 6135 17088 6408 17116
rect 6135 17085 6147 17088
rect 6089 17079 6147 17085
rect 6638 17076 6644 17128
rect 6696 17076 6702 17128
rect 2424 17020 3188 17048
rect 1854 16940 1860 16992
rect 1912 16940 1918 16992
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 2593 16983 2651 16989
rect 2593 16980 2605 16983
rect 2096 16952 2605 16980
rect 2096 16940 2102 16952
rect 2593 16949 2605 16952
rect 2639 16949 2651 16983
rect 3160 16980 3188 17020
rect 3510 17008 3516 17060
rect 3568 17008 3574 17060
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17017 3663 17051
rect 3605 17011 3663 17017
rect 3620 16980 3648 17011
rect 3694 17008 3700 17060
rect 3752 17008 3758 17060
rect 3988 17020 4476 17048
rect 3988 16992 4016 17020
rect 3160 16952 3648 16980
rect 3881 16983 3939 16989
rect 2593 16943 2651 16949
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 3970 16980 3976 16992
rect 3927 16952 3976 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4448 16980 4476 17020
rect 5718 17008 5724 17060
rect 5776 17008 5782 17060
rect 6086 16980 6092 16992
rect 4448 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16980 6150 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6144 16952 6469 16980
rect 6144 16940 6150 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 6457 16943 6515 16949
rect 7190 16940 7196 16992
rect 7248 16940 7254 16992
rect 7576 16980 7604 17156
rect 7650 17144 7656 17196
rect 7708 17144 7714 17196
rect 8018 17144 8024 17196
rect 8076 17182 8082 17196
rect 8123 17187 8181 17193
rect 8123 17182 8135 17187
rect 8076 17154 8135 17182
rect 8076 17144 8082 17154
rect 8123 17153 8135 17154
rect 8169 17153 8181 17187
rect 8220 17184 8248 17224
rect 8386 17212 8392 17264
rect 8444 17212 8450 17264
rect 9646 17224 11652 17252
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8220 17156 8677 17184
rect 8123 17147 8181 17153
rect 8665 17153 8677 17156
rect 8711 17184 8723 17187
rect 9646 17184 9674 17224
rect 8711 17156 9674 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 11054 17144 11060 17196
rect 11112 17144 11118 17196
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11624 17184 11652 17224
rect 11882 17212 11888 17264
rect 11940 17212 11946 17264
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12802 17252 12808 17264
rect 12023 17224 12808 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 15562 17212 15568 17264
rect 15620 17252 15626 17264
rect 15838 17252 15844 17264
rect 15620 17224 15844 17252
rect 15620 17212 15626 17224
rect 15838 17212 15844 17224
rect 15896 17212 15902 17264
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 22189 17255 22247 17261
rect 16080 17224 21956 17252
rect 16080 17212 16086 17224
rect 12529 17187 12587 17193
rect 11379 17156 11560 17184
rect 11624 17156 12480 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17116 7803 17119
rect 7926 17116 7932 17128
rect 7791 17088 7932 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 8021 17051 8079 17057
rect 8021 17017 8033 17051
rect 8067 17048 8079 17051
rect 8570 17048 8576 17060
rect 8067 17020 8576 17048
rect 8067 17017 8079 17020
rect 8021 17011 8079 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 9582 17008 9588 17060
rect 9640 17048 9646 17060
rect 11532 17057 11560 17156
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12452 17116 12480 17156
rect 12529 17153 12541 17187
rect 12575 17184 12587 17187
rect 12618 17184 12624 17196
rect 12575 17156 12624 17184
rect 12575 17153 12587 17156
rect 12529 17147 12587 17153
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12452 17088 12817 17116
rect 12805 17085 12817 17088
rect 12851 17116 12863 17119
rect 13814 17116 13820 17128
rect 12851 17088 13820 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 11517 17051 11575 17057
rect 9640 17020 11468 17048
rect 9640 17008 9646 17020
rect 8386 16980 8392 16992
rect 7576 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16980 8450 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8444 16952 8769 16980
rect 8444 16940 8450 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 11146 16940 11152 16992
rect 11204 16940 11210 16992
rect 11440 16980 11468 17020
rect 11517 17017 11529 17051
rect 11563 17017 11575 17051
rect 13357 17051 13415 17057
rect 13357 17048 13369 17051
rect 11517 17011 11575 17017
rect 11624 17020 13369 17048
rect 11624 16980 11652 17020
rect 13357 17017 13369 17020
rect 13403 17017 13415 17051
rect 15120 17048 15148 17147
rect 15378 17144 15384 17196
rect 15436 17144 15442 17196
rect 15470 17144 15476 17196
rect 15528 17144 15534 17196
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15804 17156 16681 17184
rect 15804 17144 15810 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19208 17156 19625 17184
rect 19208 17144 19214 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19794 17144 19800 17196
rect 19852 17144 19858 17196
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20404 17156 20637 17184
rect 20404 17144 20410 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 21315 17156 21864 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 15344 17088 16068 17116
rect 15344 17076 15350 17088
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 15120 17020 15945 17048
rect 13357 17011 13415 17017
rect 15933 17017 15945 17020
rect 15979 17017 15991 17051
rect 16040 17048 16068 17088
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16908 17088 16957 17116
rect 16908 17076 16914 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17116 20775 17119
rect 21174 17116 21180 17128
rect 20763 17088 21180 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 21634 17076 21640 17128
rect 21692 17076 21698 17128
rect 20622 17048 20628 17060
rect 16040 17020 20628 17048
rect 15933 17011 15991 17017
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 11440 16952 11652 16980
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 12434 16980 12440 16992
rect 12391 16952 12440 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 14918 16940 14924 16992
rect 14976 16940 14982 16992
rect 15289 16983 15347 16989
rect 15289 16949 15301 16983
rect 15335 16980 15347 16983
rect 15562 16980 15568 16992
rect 15335 16952 15568 16980
rect 15335 16949 15347 16952
rect 15289 16943 15347 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 16761 16983 16819 16989
rect 16761 16949 16773 16983
rect 16807 16980 16819 16983
rect 18690 16980 18696 16992
rect 16807 16952 18696 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 19610 16940 19616 16992
rect 19668 16940 19674 16992
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 21652 16980 21680 17076
rect 21836 17057 21864 17156
rect 21821 17051 21879 17057
rect 21821 17017 21833 17051
rect 21867 17017 21879 17051
rect 21928 17048 21956 17224
rect 22189 17221 22201 17255
rect 22235 17252 22247 17255
rect 22848 17252 22876 17280
rect 22235 17224 22876 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 22370 17076 22376 17128
rect 22428 17076 22434 17128
rect 23124 17048 23152 17280
rect 23584 17193 23612 17292
rect 24394 17280 24400 17292
rect 24452 17280 24458 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 25884 17320 25912 17564
rect 25363 17292 25912 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 23658 17212 23664 17264
rect 23716 17252 23722 17264
rect 23845 17255 23903 17261
rect 23845 17252 23857 17255
rect 23716 17224 23857 17252
rect 23716 17212 23722 17224
rect 23845 17221 23857 17224
rect 23891 17221 23903 17255
rect 23845 17215 23903 17221
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17184 25559 17187
rect 25547 17156 26004 17184
rect 25547 17153 25559 17156
rect 25501 17147 25559 17153
rect 25056 17116 25084 17147
rect 25682 17116 25688 17128
rect 21928 17020 23152 17048
rect 23216 17088 24716 17116
rect 25056 17088 25688 17116
rect 21821 17011 21879 17017
rect 23216 16980 23244 17088
rect 23934 17008 23940 17060
rect 23992 17048 23998 17060
rect 24121 17051 24179 17057
rect 24121 17048 24133 17051
rect 23992 17020 24133 17048
rect 23992 17008 23998 17020
rect 24121 17017 24133 17020
rect 24167 17048 24179 17051
rect 24578 17048 24584 17060
rect 24167 17020 24584 17048
rect 24167 17017 24179 17020
rect 24121 17011 24179 17017
rect 24578 17008 24584 17020
rect 24636 17008 24642 17060
rect 24688 17048 24716 17088
rect 25682 17076 25688 17088
rect 25740 17076 25746 17128
rect 25976 17060 26004 17156
rect 25225 17051 25283 17057
rect 25225 17048 25237 17051
rect 24688 17020 25237 17048
rect 25225 17017 25237 17020
rect 25271 17017 25283 17051
rect 25225 17011 25283 17017
rect 25958 17008 25964 17060
rect 26016 17008 26022 17060
rect 21652 16952 23244 16980
rect 23385 16983 23443 16989
rect 23385 16949 23397 16983
rect 23431 16980 23443 16983
rect 24026 16980 24032 16992
rect 23431 16952 24032 16980
rect 23431 16949 23443 16952
rect 23385 16943 23443 16949
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24305 16983 24363 16989
rect 24305 16949 24317 16983
rect 24351 16980 24363 16983
rect 24854 16980 24860 16992
rect 24351 16952 24860 16980
rect 24351 16949 24363 16952
rect 24305 16943 24363 16949
rect 24854 16940 24860 16952
rect 24912 16940 24918 16992
rect 1104 16890 25852 16912
rect 1104 16838 4043 16890
rect 4095 16838 4107 16890
rect 4159 16838 4171 16890
rect 4223 16838 4235 16890
rect 4287 16838 4299 16890
rect 4351 16838 10230 16890
rect 10282 16838 10294 16890
rect 10346 16838 10358 16890
rect 10410 16838 10422 16890
rect 10474 16838 10486 16890
rect 10538 16838 16417 16890
rect 16469 16838 16481 16890
rect 16533 16838 16545 16890
rect 16597 16838 16609 16890
rect 16661 16838 16673 16890
rect 16725 16838 22604 16890
rect 22656 16838 22668 16890
rect 22720 16838 22732 16890
rect 22784 16838 22796 16890
rect 22848 16838 22860 16890
rect 22912 16838 25852 16890
rect 1104 16816 25852 16838
rect 1670 16736 1676 16788
rect 1728 16736 1734 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3510 16776 3516 16788
rect 2924 16748 3516 16776
rect 2924 16736 2930 16748
rect 3510 16736 3516 16748
rect 3568 16776 3574 16788
rect 3568 16748 5304 16776
rect 3568 16736 3574 16748
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 1688 16640 1716 16736
rect 4246 16708 4252 16720
rect 3252 16680 4252 16708
rect 1627 16612 1716 16640
rect 1857 16643 1915 16649
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 3252 16640 3280 16680
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 4522 16668 4528 16720
rect 4580 16668 4586 16720
rect 5276 16717 5304 16748
rect 5994 16736 6000 16788
rect 6052 16736 6058 16788
rect 6362 16736 6368 16788
rect 6420 16736 6426 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 11054 16776 11060 16788
rect 10459 16748 11060 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11314 16779 11372 16785
rect 11314 16776 11326 16779
rect 11204 16748 11326 16776
rect 11204 16736 11210 16748
rect 11314 16745 11326 16748
rect 11360 16745 11372 16779
rect 16942 16776 16948 16788
rect 11314 16739 11372 16745
rect 13740 16748 16948 16776
rect 5261 16711 5319 16717
rect 5261 16677 5273 16711
rect 5307 16708 5319 16711
rect 5534 16708 5540 16720
rect 5307 16680 5540 16708
rect 5307 16677 5319 16680
rect 5261 16671 5319 16677
rect 5534 16668 5540 16680
rect 5592 16708 5598 16720
rect 5813 16711 5871 16717
rect 5813 16708 5825 16711
rect 5592 16680 5825 16708
rect 5592 16668 5598 16680
rect 5813 16677 5825 16680
rect 5859 16708 5871 16711
rect 10321 16711 10379 16717
rect 5859 16680 10272 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 1903 16612 3280 16640
rect 3329 16643 3387 16649
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3375 16612 3801 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 4893 16643 4951 16649
rect 3789 16603 3847 16609
rect 4356 16612 4844 16640
rect 3602 16532 3608 16584
rect 3660 16532 3666 16584
rect 3694 16532 3700 16584
rect 3752 16572 3758 16584
rect 4356 16572 4384 16612
rect 4816 16581 4844 16612
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5442 16640 5448 16652
rect 4939 16612 5448 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 9582 16640 9588 16652
rect 5828 16612 6316 16640
rect 3752 16544 4384 16572
rect 4801 16575 4859 16581
rect 3752 16532 3758 16544
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 5828 16572 5856 16612
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 4801 16535 4859 16541
rect 5368 16544 5856 16572
rect 5920 16544 6193 16572
rect 3082 16476 3188 16504
rect 3160 16436 3188 16476
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 4525 16507 4583 16513
rect 4525 16504 4537 16507
rect 3844 16476 4537 16504
rect 3844 16464 3850 16476
rect 4525 16473 4537 16476
rect 4571 16504 4583 16507
rect 4614 16504 4620 16516
rect 4571 16476 4620 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 4614 16464 4620 16476
rect 4672 16464 4678 16516
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3160 16408 3433 16436
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 5368 16445 5396 16544
rect 5442 16464 5448 16516
rect 5500 16464 5506 16516
rect 5920 16445 5948 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6288 16572 6316 16612
rect 8128 16612 9588 16640
rect 8128 16581 8156 16612
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10244 16640 10272 16680
rect 10321 16677 10333 16711
rect 10367 16708 10379 16711
rect 10594 16708 10600 16720
rect 10367 16680 10600 16708
rect 10367 16677 10379 16680
rect 10321 16671 10379 16677
rect 10594 16668 10600 16680
rect 10652 16668 10658 16720
rect 10781 16711 10839 16717
rect 10781 16677 10793 16711
rect 10827 16677 10839 16711
rect 10781 16671 10839 16677
rect 10410 16640 10416 16652
rect 10244 16612 10416 16640
rect 10410 16600 10416 16612
rect 10468 16640 10474 16652
rect 10796 16640 10824 16671
rect 10468 16612 10824 16640
rect 10468 16600 10474 16612
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 13740 16649 13768 16748
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 18064 16748 19380 16776
rect 14550 16668 14556 16720
rect 14608 16708 14614 16720
rect 16850 16708 16856 16720
rect 14608 16680 16856 16708
rect 14608 16668 14614 16680
rect 16850 16668 16856 16680
rect 16908 16708 16914 16720
rect 16908 16680 17908 16708
rect 16908 16668 16914 16680
rect 13725 16643 13783 16649
rect 13725 16640 13737 16643
rect 12124 16612 13737 16640
rect 12124 16600 12130 16612
rect 13725 16609 13737 16612
rect 13771 16609 13783 16643
rect 13725 16603 13783 16609
rect 14737 16643 14795 16649
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 14918 16640 14924 16652
rect 14783 16612 14924 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 15381 16643 15439 16649
rect 15381 16609 15393 16643
rect 15427 16640 15439 16643
rect 15562 16640 15568 16652
rect 15427 16612 15568 16640
rect 15427 16609 15439 16612
rect 15381 16603 15439 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15746 16640 15752 16652
rect 15703 16612 15752 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 17880 16649 17908 16680
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16609 17923 16643
rect 17865 16603 17923 16609
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6288 16544 6561 16572
rect 6181 16535 6239 16541
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 8297 16575 8355 16581
rect 8297 16541 8309 16575
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 8018 16464 8024 16516
rect 8076 16504 8082 16516
rect 8220 16504 8248 16535
rect 8076 16476 8248 16504
rect 8312 16504 8340 16535
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8754 16532 8760 16584
rect 8812 16532 8818 16584
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 11057 16575 11115 16581
rect 8996 16544 10548 16572
rect 8996 16532 9002 16544
rect 10520 16513 10548 16544
rect 11057 16541 11069 16575
rect 11103 16541 11115 16575
rect 11057 16535 11115 16541
rect 8665 16507 8723 16513
rect 8665 16504 8677 16507
rect 8312 16476 8677 16504
rect 8076 16464 8082 16476
rect 8665 16473 8677 16476
rect 8711 16473 8723 16507
rect 8665 16467 8723 16473
rect 9953 16507 10011 16513
rect 9953 16473 9965 16507
rect 9999 16504 10011 16507
rect 10505 16507 10563 16513
rect 9999 16476 10088 16504
rect 9999 16473 10011 16476
rect 9953 16467 10011 16473
rect 10060 16448 10088 16476
rect 10505 16473 10517 16507
rect 10551 16504 10563 16507
rect 10686 16504 10692 16516
rect 10551 16476 10692 16504
rect 10551 16473 10563 16476
rect 10505 16467 10563 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 11072 16504 11100 16535
rect 12434 16532 12440 16584
rect 12492 16532 12498 16584
rect 14642 16532 14648 16584
rect 14700 16532 14706 16584
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 11330 16504 11336 16516
rect 11072 16476 11336 16504
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 13446 16464 13452 16516
rect 13504 16504 13510 16516
rect 13541 16507 13599 16513
rect 13541 16504 13553 16507
rect 13504 16476 13553 16504
rect 13504 16464 13510 16476
rect 13541 16473 13553 16476
rect 13587 16504 13599 16507
rect 15304 16504 15332 16535
rect 16206 16532 16212 16584
rect 16264 16532 16270 16584
rect 18064 16581 18092 16748
rect 18785 16711 18843 16717
rect 18785 16677 18797 16711
rect 18831 16708 18843 16711
rect 19352 16708 19380 16748
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 19889 16779 19947 16785
rect 19889 16776 19901 16779
rect 19852 16748 19901 16776
rect 19852 16736 19858 16748
rect 19889 16745 19901 16748
rect 19935 16745 19947 16779
rect 19889 16739 19947 16745
rect 20898 16736 20904 16788
rect 20956 16736 20962 16788
rect 21729 16779 21787 16785
rect 21729 16745 21741 16779
rect 21775 16776 21787 16779
rect 21910 16776 21916 16788
rect 21775 16748 21916 16776
rect 21775 16745 21787 16748
rect 21729 16739 21787 16745
rect 19981 16711 20039 16717
rect 19981 16708 19993 16711
rect 18831 16680 19288 16708
rect 19352 16680 19993 16708
rect 18831 16677 18843 16680
rect 18785 16671 18843 16677
rect 18230 16600 18236 16652
rect 18288 16600 18294 16652
rect 18690 16600 18696 16652
rect 18748 16600 18754 16652
rect 19260 16649 19288 16680
rect 19981 16677 19993 16680
rect 20027 16677 20039 16711
rect 20916 16708 20944 16736
rect 19981 16671 20039 16677
rect 20456 16680 20944 16708
rect 20456 16649 20484 16680
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 20441 16643 20499 16649
rect 20441 16609 20453 16643
rect 20487 16609 20499 16643
rect 20441 16603 20499 16609
rect 20622 16600 20628 16652
rect 20680 16600 20686 16652
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16640 20867 16643
rect 21361 16643 21419 16649
rect 20855 16612 21312 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18196 16544 18337 16572
rect 18196 16532 18202 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18414 16532 18420 16584
rect 18472 16532 18478 16584
rect 18708 16572 18736 16600
rect 19061 16575 19119 16581
rect 19061 16572 19073 16575
rect 18708 16544 19073 16572
rect 19061 16541 19073 16544
rect 19107 16572 19119 16575
rect 19794 16572 19800 16584
rect 19107 16544 19800 16572
rect 19107 16541 19119 16544
rect 19061 16535 19119 16541
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20404 16544 21005 16572
rect 20404 16532 20410 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 21284 16572 21312 16612
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 21744 16640 21772 16739
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22097 16779 22155 16785
rect 22097 16745 22109 16779
rect 22143 16745 22155 16779
rect 22097 16739 22155 16745
rect 22112 16708 22140 16739
rect 22186 16708 22192 16720
rect 22112 16680 22192 16708
rect 22186 16668 22192 16680
rect 22244 16668 22250 16720
rect 22370 16668 22376 16720
rect 22428 16708 22434 16720
rect 22465 16711 22523 16717
rect 22465 16708 22477 16711
rect 22428 16680 22477 16708
rect 22428 16668 22434 16680
rect 22465 16677 22477 16680
rect 22511 16677 22523 16711
rect 22465 16671 22523 16677
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 24670 16708 24676 16720
rect 23716 16680 24676 16708
rect 23716 16668 23722 16680
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 23842 16640 23848 16652
rect 21407 16612 21772 16640
rect 23676 16612 23848 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 21284 16544 21465 16572
rect 20993 16535 21051 16541
rect 21453 16541 21465 16544
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 15378 16504 15384 16516
rect 13587 16476 15240 16504
rect 15304 16476 15384 16504
rect 13587 16473 13599 16476
rect 13541 16467 13599 16473
rect 4433 16439 4491 16445
rect 4433 16436 4445 16439
rect 4120 16408 4445 16436
rect 4120 16396 4126 16408
rect 4433 16405 4445 16408
rect 4479 16436 4491 16439
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4479 16408 4721 16436
rect 4479 16405 4491 16408
rect 4433 16399 4491 16405
rect 4709 16405 4721 16408
rect 4755 16405 4767 16439
rect 4709 16399 4767 16405
rect 5353 16439 5411 16445
rect 5353 16405 5365 16439
rect 5399 16405 5411 16439
rect 5353 16399 5411 16405
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16405 5963 16439
rect 5905 16399 5963 16405
rect 7834 16396 7840 16448
rect 7892 16396 7898 16448
rect 10042 16396 10048 16448
rect 10100 16396 10106 16448
rect 10965 16439 11023 16445
rect 10965 16405 10977 16439
rect 11011 16436 11023 16439
rect 12618 16436 12624 16448
rect 11011 16408 12624 16436
rect 11011 16405 11023 16408
rect 10965 16399 11023 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12802 16396 12808 16448
rect 12860 16396 12866 16448
rect 13170 16396 13176 16448
rect 13228 16396 13234 16448
rect 13633 16439 13691 16445
rect 13633 16405 13645 16439
rect 13679 16436 13691 16439
rect 14182 16436 14188 16448
rect 13679 16408 14188 16436
rect 13679 16405 13691 16408
rect 13633 16399 13691 16405
rect 14182 16396 14188 16408
rect 14240 16396 14246 16448
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 15212 16436 15240 16476
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 16761 16507 16819 16513
rect 16761 16473 16773 16507
rect 16807 16504 16819 16507
rect 18785 16507 18843 16513
rect 16807 16476 17908 16504
rect 16807 16473 16819 16476
rect 16761 16467 16819 16473
rect 17770 16436 17776 16448
rect 15212 16408 17776 16436
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 17880 16436 17908 16476
rect 18785 16473 18797 16507
rect 18831 16504 18843 16507
rect 19426 16504 19432 16516
rect 18831 16476 19432 16504
rect 18831 16473 18843 16476
rect 18785 16467 18843 16473
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 21468 16504 21496 16535
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 21994 16577 22052 16583
rect 21994 16574 22006 16577
rect 21928 16572 22006 16574
rect 21876 16546 22006 16572
rect 21876 16544 21956 16546
rect 21876 16532 21882 16544
rect 21994 16543 22006 16546
rect 22040 16543 22052 16577
rect 23676 16572 23704 16612
rect 23842 16600 23848 16612
rect 23900 16600 23906 16652
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24946 16640 24952 16652
rect 24535 16612 24952 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 21994 16537 22052 16543
rect 22388 16544 23704 16572
rect 23753 16575 23811 16581
rect 22278 16504 22284 16516
rect 19536 16476 21036 16504
rect 21468 16476 22284 16504
rect 18969 16439 19027 16445
rect 18969 16436 18981 16439
rect 17880 16408 18981 16436
rect 18969 16405 18981 16408
rect 19015 16405 19027 16439
rect 18969 16399 19027 16405
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 19536 16436 19564 16476
rect 19116 16408 19564 16436
rect 20349 16439 20407 16445
rect 19116 16396 19122 16408
rect 20349 16405 20361 16439
rect 20395 16436 20407 16439
rect 20898 16436 20904 16448
rect 20395 16408 20904 16436
rect 20395 16405 20407 16408
rect 20349 16399 20407 16405
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 21008 16445 21036 16476
rect 22278 16464 22284 16476
rect 22336 16464 22342 16516
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16405 21051 16439
rect 20993 16399 21051 16405
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 21913 16439 21971 16445
rect 21913 16436 21925 16439
rect 21232 16408 21925 16436
rect 21232 16396 21238 16408
rect 21913 16405 21925 16408
rect 21959 16405 21971 16439
rect 21913 16399 21971 16405
rect 22002 16396 22008 16448
rect 22060 16436 22066 16448
rect 22388 16436 22416 16544
rect 23753 16541 23765 16575
rect 23799 16572 23811 16575
rect 23934 16572 23940 16584
rect 23799 16544 23940 16572
rect 23799 16541 23811 16544
rect 23753 16535 23811 16541
rect 23934 16532 23940 16544
rect 23992 16532 23998 16584
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16541 24087 16575
rect 24029 16535 24087 16541
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 24044 16504 24072 16535
rect 24854 16532 24860 16584
rect 24912 16572 24918 16584
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 24912 16544 25329 16572
rect 24912 16532 24918 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 22888 16476 24072 16504
rect 22888 16464 22894 16476
rect 22060 16408 22416 16436
rect 22060 16396 22066 16408
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 23569 16439 23627 16445
rect 23569 16436 23581 16439
rect 22520 16408 23581 16436
rect 22520 16396 22526 16408
rect 23569 16405 23581 16408
rect 23615 16405 23627 16439
rect 23569 16399 23627 16405
rect 23842 16396 23848 16448
rect 23900 16396 23906 16448
rect 25038 16396 25044 16448
rect 25096 16396 25102 16448
rect 25133 16439 25191 16445
rect 25133 16405 25145 16439
rect 25179 16436 25191 16439
rect 25222 16436 25228 16448
rect 25179 16408 25228 16436
rect 25179 16405 25191 16408
rect 25133 16399 25191 16405
rect 25222 16396 25228 16408
rect 25280 16396 25286 16448
rect 1104 16346 25852 16368
rect 1104 16294 4703 16346
rect 4755 16294 4767 16346
rect 4819 16294 4831 16346
rect 4883 16294 4895 16346
rect 4947 16294 4959 16346
rect 5011 16294 10890 16346
rect 10942 16294 10954 16346
rect 11006 16294 11018 16346
rect 11070 16294 11082 16346
rect 11134 16294 11146 16346
rect 11198 16294 17077 16346
rect 17129 16294 17141 16346
rect 17193 16294 17205 16346
rect 17257 16294 17269 16346
rect 17321 16294 17333 16346
rect 17385 16294 23264 16346
rect 23316 16294 23328 16346
rect 23380 16294 23392 16346
rect 23444 16294 23456 16346
rect 23508 16294 23520 16346
rect 23572 16294 25852 16346
rect 1104 16272 25852 16294
rect 3053 16235 3111 16241
rect 3053 16201 3065 16235
rect 3099 16232 3111 16235
rect 3602 16232 3608 16244
rect 3099 16204 3608 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 3602 16192 3608 16204
rect 3660 16192 3666 16244
rect 4246 16192 4252 16244
rect 4304 16192 4310 16244
rect 4522 16192 4528 16244
rect 4580 16192 4586 16244
rect 7834 16192 7840 16244
rect 7892 16192 7898 16244
rect 8018 16192 8024 16244
rect 8076 16232 8082 16244
rect 8570 16232 8576 16244
rect 8076 16204 8576 16232
rect 8076 16192 8082 16204
rect 8570 16192 8576 16204
rect 8628 16232 8634 16244
rect 9214 16232 9220 16244
rect 8628 16204 9220 16232
rect 8628 16192 8634 16204
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9677 16235 9735 16241
rect 9677 16232 9689 16235
rect 9548 16204 9689 16232
rect 9548 16192 9554 16204
rect 9677 16201 9689 16204
rect 9723 16201 9735 16235
rect 9677 16195 9735 16201
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10778 16232 10784 16244
rect 10459 16204 10784 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11020 16204 11560 16232
rect 11020 16192 11026 16204
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 3145 16167 3203 16173
rect 3145 16164 3157 16167
rect 2832 16136 3157 16164
rect 2832 16124 2838 16136
rect 3145 16133 3157 16136
rect 3191 16133 3203 16167
rect 3145 16127 3203 16133
rect 3329 16167 3387 16173
rect 3329 16133 3341 16167
rect 3375 16164 3387 16167
rect 4062 16164 4068 16176
rect 3375 16136 4068 16164
rect 3375 16133 3387 16136
rect 3329 16127 3387 16133
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 4540 16164 4568 16192
rect 4172 16136 4568 16164
rect 4172 16105 4200 16136
rect 4614 16124 4620 16176
rect 4672 16124 4678 16176
rect 7852 16164 7880 16192
rect 11532 16176 11560 16204
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 12253 16235 12311 16241
rect 12253 16232 12265 16235
rect 11756 16204 12265 16232
rect 11756 16192 11762 16204
rect 12253 16201 12265 16204
rect 12299 16201 12311 16235
rect 12253 16195 12311 16201
rect 15746 16192 15752 16244
rect 15804 16192 15810 16244
rect 17494 16232 17500 16244
rect 16040 16204 17500 16232
rect 8205 16167 8263 16173
rect 8205 16164 8217 16167
rect 7852 16136 8217 16164
rect 8205 16133 8217 16136
rect 8251 16133 8263 16167
rect 11422 16164 11428 16176
rect 8205 16127 8263 16133
rect 9646 16136 11428 16164
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 4157 16099 4215 16105
rect 1535 16068 2268 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 2240 15901 2268 16068
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 2498 15988 2504 16040
rect 2556 16028 2562 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2556 16000 2605 16028
rect 2556 15988 2562 16000
rect 2593 15997 2605 16000
rect 2639 16028 2651 16031
rect 2639 16000 3004 16028
rect 2639 15997 2651 16000
rect 2593 15991 2651 15997
rect 2866 15920 2872 15972
rect 2924 15920 2930 15972
rect 2976 15960 3004 16000
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3513 16031 3571 16037
rect 3513 16028 3525 16031
rect 3108 16000 3525 16028
rect 3108 15988 3114 16000
rect 3513 15997 3525 16000
rect 3559 16028 3571 16031
rect 4356 16028 4384 16059
rect 3559 16000 4384 16028
rect 4632 16028 4660 16124
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 6972 16068 7941 16096
rect 6972 16056 6978 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9646 16028 9674 16136
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 11514 16124 11520 16176
rect 11572 16124 11578 16176
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 11940 16136 12112 16164
rect 11940 16124 11946 16136
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 11054 16096 11060 16108
rect 10560 16068 11060 16096
rect 10560 16056 10566 16068
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11790 16056 11796 16108
rect 11848 16056 11854 16108
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 12084 16105 12112 16136
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 12676 16136 13202 16164
rect 12676 16124 12682 16136
rect 15470 16124 15476 16176
rect 15528 16164 15534 16176
rect 15657 16167 15715 16173
rect 15657 16164 15669 16167
rect 15528 16136 15669 16164
rect 15528 16124 15534 16136
rect 15657 16133 15669 16136
rect 15703 16164 15715 16167
rect 16040 16164 16068 16204
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17770 16192 17776 16244
rect 17828 16232 17834 16244
rect 17828 16204 18828 16232
rect 17828 16192 17834 16204
rect 15703 16136 16068 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 16206 16124 16212 16176
rect 16264 16124 16270 16176
rect 17586 16164 17592 16176
rect 17144 16136 17592 16164
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16065 12127 16099
rect 16224 16096 16252 16124
rect 17144 16105 17172 16136
rect 17586 16124 17592 16136
rect 17644 16124 17650 16176
rect 18230 16124 18236 16176
rect 18288 16124 18294 16176
rect 18800 16164 18828 16204
rect 18966 16192 18972 16244
rect 19024 16192 19030 16244
rect 19613 16235 19671 16241
rect 19613 16201 19625 16235
rect 19659 16232 19671 16235
rect 20346 16232 20352 16244
rect 19659 16204 20352 16232
rect 19659 16201 19671 16204
rect 19613 16195 19671 16201
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 22002 16232 22008 16244
rect 20456 16204 22008 16232
rect 20456 16164 20484 16204
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 22281 16235 22339 16241
rect 22281 16232 22293 16235
rect 22204 16204 22293 16232
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 18800 16136 20484 16164
rect 20548 16136 21097 16164
rect 12069 16059 12127 16065
rect 13924 16068 16252 16096
rect 17129 16099 17187 16105
rect 4632 16000 9674 16028
rect 9953 16031 10011 16037
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 9999 16000 10088 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 3142 15960 3148 15972
rect 2976 15932 3148 15960
rect 3142 15920 3148 15932
rect 3200 15920 3206 15972
rect 10060 15904 10088 16000
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10468 16000 10824 16028
rect 10468 15988 10474 16000
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 10594 15960 10600 15972
rect 10367 15932 10600 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 10594 15920 10600 15932
rect 10652 15920 10658 15972
rect 10796 15960 10824 16000
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11992 16000 12449 16028
rect 11146 15960 11152 15972
rect 10796 15932 11152 15960
rect 11146 15920 11152 15932
rect 11204 15920 11210 15972
rect 11348 15960 11376 15988
rect 11992 15960 12020 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12710 15988 12716 16040
rect 12768 15988 12774 16040
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13924 16028 13952 16068
rect 17129 16065 17141 16099
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 19153 16099 19211 16105
rect 19153 16065 19165 16099
rect 19199 16096 19211 16099
rect 19334 16096 19340 16108
rect 19199 16068 19340 16096
rect 19199 16065 19211 16068
rect 19153 16059 19211 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19610 16056 19616 16108
rect 19668 16096 19674 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19668 16068 19717 16096
rect 19668 16056 19674 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 20548 16096 20576 16136
rect 21085 16133 21097 16136
rect 21131 16133 21143 16167
rect 21085 16127 21143 16133
rect 21818 16124 21824 16176
rect 21876 16124 21882 16176
rect 19852 16068 20576 16096
rect 20993 16099 21051 16105
rect 19852 16056 19858 16068
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21039 16068 21588 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 12860 16000 13952 16028
rect 12860 15988 12866 16000
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15746 16028 15752 16040
rect 15344 16000 15752 16028
rect 15344 15988 15350 16000
rect 15746 15988 15752 16000
rect 15804 16028 15810 16040
rect 15841 16031 15899 16037
rect 15841 16028 15853 16031
rect 15804 16000 15853 16028
rect 15804 15988 15810 16000
rect 15841 15997 15853 16000
rect 15887 15997 15899 16031
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 15841 15991 15899 15997
rect 15948 16000 17233 16028
rect 11348 15932 12020 15960
rect 12084 15932 12434 15960
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 5626 15892 5632 15904
rect 2271 15864 5632 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5718 15852 5724 15904
rect 5776 15852 5782 15904
rect 10042 15852 10048 15904
rect 10100 15852 10106 15904
rect 10612 15892 10640 15920
rect 10689 15895 10747 15901
rect 10689 15892 10701 15895
rect 10612 15864 10701 15892
rect 10689 15861 10701 15864
rect 10735 15861 10747 15895
rect 10689 15855 10747 15861
rect 11330 15852 11336 15904
rect 11388 15852 11394 15904
rect 12084 15901 12112 15932
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15861 12127 15895
rect 12406 15892 12434 15932
rect 15948 15904 15976 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17221 15991 17279 15997
rect 17328 16000 17509 16028
rect 16945 15963 17003 15969
rect 16945 15929 16957 15963
rect 16991 15960 17003 15963
rect 17328 15960 17356 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 18138 16028 18144 16040
rect 17644 16000 18144 16028
rect 17644 15988 17650 16000
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 21082 16028 21088 16040
rect 18840 16000 21088 16028
rect 18840 15988 18846 16000
rect 21082 15988 21088 16000
rect 21140 16028 21146 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 21140 16000 21189 16028
rect 21140 15988 21146 16000
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 16991 15932 17356 15960
rect 16991 15929 17003 15932
rect 16945 15923 17003 15929
rect 18506 15920 18512 15972
rect 18564 15960 18570 15972
rect 19610 15960 19616 15972
rect 18564 15932 19616 15960
rect 18564 15920 18570 15932
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 13446 15892 13452 15904
rect 12406 15864 13452 15892
rect 12069 15855 12127 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 14182 15852 14188 15904
rect 14240 15852 14246 15904
rect 15286 15852 15292 15904
rect 15344 15852 15350 15904
rect 15930 15852 15936 15904
rect 15988 15852 15994 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 19334 15892 19340 15904
rect 16264 15864 19340 15892
rect 16264 15852 16270 15864
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19426 15852 19432 15904
rect 19484 15852 19490 15904
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 19944 15864 20361 15892
rect 19944 15852 19950 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20349 15855 20407 15861
rect 20625 15895 20683 15901
rect 20625 15861 20637 15895
rect 20671 15892 20683 15895
rect 20714 15892 20720 15904
rect 20671 15864 20720 15892
rect 20671 15861 20683 15864
rect 20625 15855 20683 15861
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 21560 15892 21588 16068
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22204 16096 22232 16204
rect 22281 16201 22293 16204
rect 22327 16201 22339 16235
rect 22281 16195 22339 16201
rect 22830 16192 22836 16244
rect 22888 16192 22894 16244
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 23382 16232 23388 16244
rect 23339 16204 23388 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23842 16192 23848 16244
rect 23900 16192 23906 16244
rect 25409 16235 25467 16241
rect 25409 16201 25421 16235
rect 25455 16232 25467 16235
rect 26142 16232 26148 16244
rect 25455 16204 26148 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 23860 16164 23888 16192
rect 23937 16167 23995 16173
rect 23937 16164 23949 16167
rect 23860 16136 23949 16164
rect 23937 16133 23949 16136
rect 23983 16133 23995 16167
rect 25222 16164 25228 16176
rect 25162 16136 25228 16164
rect 23937 16127 23995 16133
rect 25222 16124 25228 16136
rect 25280 16124 25286 16176
rect 21968 16068 22232 16096
rect 21968 16056 21974 16068
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 23382 16028 23388 16040
rect 22152 16000 23388 16028
rect 22152 15988 22158 16000
rect 23382 15988 23388 16000
rect 23440 15988 23446 16040
rect 23661 16031 23719 16037
rect 23661 15997 23673 16031
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 22186 15920 22192 15972
rect 22244 15920 22250 15972
rect 22278 15920 22284 15972
rect 22336 15960 22342 15972
rect 23014 15960 23020 15972
rect 22336 15932 23020 15960
rect 22336 15920 22342 15932
rect 23014 15920 23020 15932
rect 23072 15960 23078 15972
rect 23676 15960 23704 15991
rect 25222 15988 25228 16040
rect 25280 16028 25286 16040
rect 25424 16028 25452 16195
rect 26142 16192 26148 16204
rect 26200 16192 26206 16244
rect 25280 16000 25452 16028
rect 25280 15988 25286 16000
rect 23072 15932 23704 15960
rect 23072 15920 23078 15932
rect 25498 15892 25504 15904
rect 21560 15864 25504 15892
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 1104 15802 25852 15824
rect 1104 15750 4043 15802
rect 4095 15750 4107 15802
rect 4159 15750 4171 15802
rect 4223 15750 4235 15802
rect 4287 15750 4299 15802
rect 4351 15750 10230 15802
rect 10282 15750 10294 15802
rect 10346 15750 10358 15802
rect 10410 15750 10422 15802
rect 10474 15750 10486 15802
rect 10538 15750 16417 15802
rect 16469 15750 16481 15802
rect 16533 15750 16545 15802
rect 16597 15750 16609 15802
rect 16661 15750 16673 15802
rect 16725 15750 22604 15802
rect 22656 15750 22668 15802
rect 22720 15750 22732 15802
rect 22784 15750 22796 15802
rect 22848 15750 22860 15802
rect 22912 15750 25852 15802
rect 1104 15728 25852 15750
rect 6914 15688 6920 15700
rect 5000 15660 6920 15688
rect 3786 15620 3792 15632
rect 2700 15592 3792 15620
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2700 15493 2728 15592
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 2884 15524 3372 15552
rect 2884 15493 2912 15524
rect 3344 15496 3372 15524
rect 3510 15512 3516 15564
rect 3568 15552 3574 15564
rect 5000 15561 5028 15660
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 9364 15660 9413 15688
rect 9364 15648 9370 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 9401 15651 9459 15657
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 9950 15688 9956 15700
rect 9640 15660 9956 15688
rect 9640 15648 9646 15660
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 10928 15660 11621 15688
rect 10928 15648 10934 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 12618 15688 12624 15700
rect 12575 15660 12624 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12768 15660 12909 15688
rect 12768 15648 12774 15660
rect 12897 15657 12909 15660
rect 12943 15657 12955 15691
rect 19058 15688 19064 15700
rect 12897 15651 12955 15657
rect 16040 15660 19064 15688
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 16040 15620 16068 15660
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 19508 15691 19566 15697
rect 19508 15657 19520 15691
rect 19554 15688 19566 15691
rect 19886 15688 19892 15700
rect 19554 15660 19892 15688
rect 19554 15657 19566 15660
rect 19508 15651 19566 15657
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 20993 15691 21051 15697
rect 20993 15688 21005 15691
rect 20956 15660 21005 15688
rect 20956 15648 20962 15660
rect 20993 15657 21005 15660
rect 21039 15688 21051 15691
rect 22186 15688 22192 15700
rect 21039 15660 22192 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 22388 15660 22600 15688
rect 7984 15592 16068 15620
rect 7984 15580 7990 15592
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 18874 15620 18880 15632
rect 17552 15592 18880 15620
rect 17552 15580 17558 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 22388 15620 22416 15660
rect 22204 15592 22416 15620
rect 4985 15555 5043 15561
rect 3568 15524 4844 15552
rect 3568 15512 3574 15524
rect 2685 15487 2743 15493
rect 2685 15484 2697 15487
rect 2096 15456 2697 15484
rect 2096 15444 2102 15456
rect 2685 15453 2697 15456
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3050 15484 3056 15496
rect 3007 15456 3056 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 3252 15416 3280 15447
rect 3326 15444 3332 15496
rect 3384 15484 3390 15496
rect 4816 15493 4844 15524
rect 4985 15521 4997 15555
rect 5031 15521 5043 15555
rect 4985 15515 5043 15521
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 11238 15552 11244 15564
rect 5684 15524 11244 15552
rect 5684 15512 5690 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11388 15524 12434 15552
rect 11388 15512 11394 15524
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3384 15456 3801 15484
rect 3384 15444 3390 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 8202 15484 8208 15496
rect 7055 15456 8208 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 4433 15419 4491 15425
rect 4433 15416 4445 15419
rect 3252 15388 4445 15416
rect 4433 15385 4445 15388
rect 4479 15385 4491 15419
rect 4433 15379 4491 15385
rect 2501 15351 2559 15357
rect 2501 15317 2513 15351
rect 2547 15348 2559 15351
rect 2774 15348 2780 15360
rect 2547 15320 2780 15348
rect 2547 15317 2559 15320
rect 2501 15311 2559 15317
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 3145 15351 3203 15357
rect 3145 15317 3157 15351
rect 3191 15348 3203 15351
rect 3510 15348 3516 15360
rect 3191 15320 3516 15348
rect 3191 15317 3203 15320
rect 3145 15311 3203 15317
rect 3510 15308 3516 15320
rect 3568 15348 3574 15360
rect 4632 15348 4660 15447
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 9122 15484 9128 15496
rect 8536 15456 9128 15484
rect 8536 15444 8542 15456
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 9950 15484 9956 15496
rect 9631 15456 9956 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10962 15484 10968 15496
rect 10367 15456 10968 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 11606 15484 11612 15496
rect 11471 15456 11612 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 12406 15484 12434 15524
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14608 15524 14933 15552
rect 14608 15512 14614 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15286 15512 15292 15564
rect 15344 15512 15350 15564
rect 15930 15512 15936 15564
rect 15988 15552 15994 15564
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 15988 15524 19257 15552
rect 15988 15512 15994 15524
rect 19245 15521 19257 15524
rect 19291 15552 19303 15555
rect 19291 15524 21312 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12406 15456 12725 15484
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13188 15484 13216 15512
rect 13127 15456 13216 15484
rect 15105 15487 15163 15493
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 15105 15453 15117 15487
rect 15151 15484 15163 15487
rect 15304 15484 15332 15512
rect 15151 15456 15332 15484
rect 15151 15453 15163 15456
rect 15105 15447 15163 15453
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18104 15456 18705 15484
rect 18104 15444 18110 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 4709 15419 4767 15425
rect 4709 15385 4721 15419
rect 4755 15416 4767 15419
rect 5261 15419 5319 15425
rect 5261 15416 5273 15419
rect 4755 15388 5273 15416
rect 4755 15385 4767 15388
rect 4709 15379 4767 15385
rect 5261 15385 5273 15388
rect 5307 15385 5319 15419
rect 5261 15379 5319 15385
rect 5718 15376 5724 15428
rect 5776 15376 5782 15428
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 16209 15419 16267 15425
rect 16209 15416 16221 15419
rect 16172 15388 16221 15416
rect 16172 15376 16178 15388
rect 16209 15385 16221 15388
rect 16255 15385 16267 15419
rect 16209 15379 16267 15385
rect 16298 15376 16304 15428
rect 16356 15416 16362 15428
rect 16356 15388 16698 15416
rect 16356 15376 16362 15388
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 17957 15419 18015 15425
rect 17957 15416 17969 15419
rect 17644 15388 17969 15416
rect 17644 15376 17650 15388
rect 17957 15385 17969 15388
rect 18003 15385 18015 15419
rect 17957 15379 18015 15385
rect 18325 15419 18383 15425
rect 18325 15385 18337 15419
rect 18371 15416 18383 15419
rect 18782 15416 18788 15428
rect 18371 15388 18788 15416
rect 18371 15385 18383 15388
rect 18325 15379 18383 15385
rect 3568 15320 4660 15348
rect 3568 15308 3574 15320
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 10042 15348 10048 15360
rect 7064 15320 10048 15348
rect 7064 15308 7070 15320
rect 10042 15308 10048 15320
rect 10100 15348 10106 15360
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10100 15320 10517 15348
rect 10100 15308 10106 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 11204 15320 11253 15348
rect 11204 15308 11210 15320
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15378 15348 15384 15360
rect 15335 15320 15384 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 18340 15348 18368 15379
rect 18782 15376 18788 15388
rect 18840 15376 18846 15428
rect 19794 15376 19800 15428
rect 19852 15416 19858 15428
rect 21284 15416 21312 15524
rect 22204 15484 22232 15592
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 22465 15555 22523 15561
rect 22465 15552 22477 15555
rect 22336 15524 22477 15552
rect 22336 15512 22342 15524
rect 22465 15521 22477 15524
rect 22511 15521 22523 15555
rect 22572 15552 22600 15660
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23440 15660 23888 15688
rect 23440 15648 23446 15660
rect 23860 15620 23888 15660
rect 23934 15648 23940 15700
rect 23992 15688 23998 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 23992 15660 24409 15688
rect 23992 15648 23998 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 24397 15651 24455 15657
rect 25406 15648 25412 15700
rect 25464 15648 25470 15700
rect 23860 15592 24992 15620
rect 23750 15552 23756 15564
rect 22572 15524 23756 15552
rect 22465 15515 22523 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24394 15552 24400 15564
rect 23992 15524 24400 15552
rect 23992 15512 23998 15524
rect 24394 15512 24400 15524
rect 24452 15552 24458 15564
rect 24964 15561 24992 15592
rect 24857 15555 24915 15561
rect 24857 15552 24869 15555
rect 24452 15524 24869 15552
rect 24452 15512 24458 15524
rect 24857 15521 24869 15524
rect 24903 15521 24915 15555
rect 24857 15515 24915 15521
rect 24949 15555 25007 15561
rect 24949 15521 24961 15555
rect 24995 15521 25007 15555
rect 24949 15515 25007 15521
rect 22373 15487 22431 15493
rect 22373 15484 22385 15487
rect 22204 15456 22385 15484
rect 22373 15453 22385 15456
rect 22419 15453 22431 15487
rect 22373 15447 22431 15453
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24544 15456 25237 15484
rect 24544 15444 24550 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 26234 15444 26240 15496
rect 26292 15444 26298 15496
rect 22278 15416 22284 15428
rect 19852 15388 20010 15416
rect 21284 15388 22284 15416
rect 19852 15376 19858 15388
rect 22278 15376 22284 15388
rect 22336 15376 22342 15428
rect 22462 15376 22468 15428
rect 22520 15416 22526 15428
rect 22741 15419 22799 15425
rect 22741 15416 22753 15419
rect 22520 15388 22753 15416
rect 22520 15376 22526 15388
rect 22741 15385 22753 15388
rect 22787 15385 22799 15419
rect 24765 15419 24823 15425
rect 22741 15379 22799 15385
rect 22848 15388 23230 15416
rect 17000 15320 18368 15348
rect 17000 15308 17006 15320
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 22002 15348 22008 15360
rect 18932 15320 22008 15348
rect 18932 15308 18938 15320
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15348 22247 15351
rect 22848 15348 22876 15388
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 26252 15416 26280 15444
rect 24811 15388 26280 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 22235 15320 22876 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 24210 15308 24216 15360
rect 24268 15308 24274 15360
rect 1104 15258 25852 15280
rect 1104 15206 4703 15258
rect 4755 15206 4767 15258
rect 4819 15206 4831 15258
rect 4883 15206 4895 15258
rect 4947 15206 4959 15258
rect 5011 15206 10890 15258
rect 10942 15206 10954 15258
rect 11006 15206 11018 15258
rect 11070 15206 11082 15258
rect 11134 15206 11146 15258
rect 11198 15206 17077 15258
rect 17129 15206 17141 15258
rect 17193 15206 17205 15258
rect 17257 15206 17269 15258
rect 17321 15206 17333 15258
rect 17385 15206 23264 15258
rect 23316 15206 23328 15258
rect 23380 15206 23392 15258
rect 23444 15206 23456 15258
rect 23508 15206 23520 15258
rect 23572 15206 25852 15258
rect 1104 15184 25852 15206
rect 1670 15104 1676 15156
rect 1728 15104 1734 15156
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 5721 15147 5779 15153
rect 2832 15116 3464 15144
rect 2832 15104 2838 15116
rect 1688 15076 1716 15104
rect 3436 15085 3464 15116
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5902 15144 5908 15156
rect 5767 15116 5908 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 9950 15104 9956 15156
rect 10008 15104 10014 15156
rect 17402 15144 17408 15156
rect 14384 15116 17408 15144
rect 1596 15048 1716 15076
rect 3421 15079 3479 15085
rect 1596 15017 1624 15048
rect 3421 15045 3433 15079
rect 3467 15045 3479 15079
rect 3421 15039 3479 15045
rect 3510 15036 3516 15088
rect 3568 15076 3574 15088
rect 3605 15079 3663 15085
rect 3605 15076 3617 15079
rect 3568 15048 3617 15076
rect 3568 15036 3574 15048
rect 3605 15045 3617 15048
rect 3651 15045 3663 15079
rect 3605 15039 3663 15045
rect 3878 15036 3884 15088
rect 3936 15076 3942 15088
rect 13081 15079 13139 15085
rect 13081 15076 13093 15079
rect 3936 15048 13093 15076
rect 3936 15036 3942 15048
rect 13081 15045 13093 15048
rect 13127 15045 13139 15079
rect 13081 15039 13139 15045
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 2958 14968 2964 15020
rect 3016 14968 3022 15020
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3200 14980 4169 15008
rect 3200 14968 3206 14980
rect 4157 14977 4169 14980
rect 4203 15008 4215 15011
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 4203 14980 5273 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 5261 14977 5273 14980
rect 5307 15008 5319 15011
rect 5442 15008 5448 15020
rect 5307 14980 5448 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 7193 15011 7251 15017
rect 6595 14980 6868 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 1854 14900 1860 14952
rect 1912 14900 1918 14952
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 2884 14912 3801 14940
rect 2406 14764 2412 14816
rect 2464 14804 2470 14816
rect 2884 14804 2912 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3326 14832 3332 14884
rect 3384 14832 3390 14884
rect 4525 14875 4583 14881
rect 4525 14841 4537 14875
rect 4571 14872 4583 14875
rect 5534 14872 5540 14884
rect 4571 14844 5540 14872
rect 4571 14841 4583 14844
rect 4525 14835 4583 14841
rect 5534 14832 5540 14844
rect 5592 14832 5598 14884
rect 6840 14881 6868 14980
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7650 15008 7656 15020
rect 7239 14980 7656 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7650 14968 7656 14980
rect 7708 15008 7714 15020
rect 11701 15011 11759 15017
rect 7708 14980 11192 15008
rect 7708 14968 7714 14980
rect 7282 14900 7288 14952
rect 7340 14900 7346 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 8478 14940 8484 14952
rect 7515 14912 8484 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 9539 14912 9674 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 6825 14875 6883 14881
rect 6825 14841 6837 14875
rect 6871 14841 6883 14875
rect 6825 14835 6883 14841
rect 2464 14776 2912 14804
rect 2464 14764 2470 14776
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5626 14804 5632 14816
rect 5132 14776 5632 14804
rect 5132 14764 5138 14776
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 6362 14764 6368 14816
rect 6420 14764 6426 14816
rect 9646 14804 9674 14912
rect 10778 14900 10784 14952
rect 10836 14900 10842 14952
rect 9861 14875 9919 14881
rect 9861 14841 9873 14875
rect 9907 14872 9919 14875
rect 10686 14872 10692 14884
rect 9907 14844 10692 14872
rect 9907 14841 9919 14844
rect 9861 14835 9919 14841
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 11054 14832 11060 14884
rect 11112 14832 11118 14884
rect 11164 14872 11192 14980
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11716 14940 11744 14971
rect 11287 14912 11744 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11164 14844 11652 14872
rect 11238 14804 11244 14816
rect 9646 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11514 14764 11520 14816
rect 11572 14764 11578 14816
rect 11624 14804 11652 14844
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 14384 14881 14412 15116
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 18230 15104 18236 15156
rect 18288 15104 18294 15156
rect 19150 15104 19156 15156
rect 19208 15104 19214 15156
rect 19794 15104 19800 15156
rect 19852 15104 19858 15156
rect 20714 15104 20720 15156
rect 20772 15104 20778 15156
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22428 15116 22937 15144
rect 22428 15104 22434 15116
rect 22925 15113 22937 15116
rect 22971 15144 22983 15147
rect 24210 15144 24216 15156
rect 22971 15116 24216 15144
rect 22971 15113 22983 15116
rect 22925 15107 22983 15113
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 24857 15147 24915 15153
rect 24857 15113 24869 15147
rect 24903 15144 24915 15147
rect 24946 15144 24952 15156
rect 24903 15116 24952 15144
rect 24903 15113 24915 15116
rect 24857 15107 24915 15113
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 15010 15036 15016 15088
rect 15068 15036 15074 15088
rect 15194 15076 15200 15088
rect 15120 15048 15200 15076
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15028 15008 15056 15036
rect 15120 15017 15148 15048
rect 15194 15036 15200 15048
rect 15252 15076 15258 15088
rect 16206 15076 16212 15088
rect 15252 15048 16212 15076
rect 15252 15036 15258 15048
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 18877 15079 18935 15085
rect 18064 15048 18644 15076
rect 18064 15020 18092 15048
rect 15378 15017 15384 15020
rect 14967 14980 15056 15008
rect 15105 15011 15163 15017
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15357 15011 15384 15017
rect 15357 14977 15369 15011
rect 15357 14971 15384 14977
rect 15378 14968 15384 14971
rect 15436 14968 15442 15020
rect 17954 15008 17960 15020
rect 16316 14980 17960 15008
rect 14734 14900 14740 14952
rect 14792 14940 14798 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 14792 14912 15025 14940
rect 14792 14900 14798 14912
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 15470 14940 15476 14952
rect 15013 14903 15071 14909
rect 15212 14912 15476 14940
rect 15212 14881 15240 14912
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 14369 14875 14427 14881
rect 14369 14872 14381 14875
rect 13596 14844 14381 14872
rect 13596 14832 13602 14844
rect 14369 14841 14381 14844
rect 14415 14841 14427 14875
rect 14369 14835 14427 14841
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14841 15255 14875
rect 15197 14835 15255 14841
rect 16316 14804 16344 14980
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18046 14968 18052 15020
rect 18104 14968 18110 15020
rect 18616 15017 18644 15048
rect 18877 15045 18889 15079
rect 18923 15076 18935 15079
rect 20254 15076 20260 15088
rect 18923 15048 20260 15076
rect 18923 15045 18935 15048
rect 18877 15039 18935 15045
rect 20254 15036 20260 15048
rect 20312 15036 20318 15088
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 17681 14943 17739 14949
rect 17681 14909 17693 14943
rect 17727 14940 17739 14943
rect 18141 14943 18199 14949
rect 17727 14912 18000 14940
rect 17727 14909 17739 14912
rect 17681 14903 17739 14909
rect 11624 14776 16344 14804
rect 17972 14804 18000 14912
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18432 14940 18460 14971
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19484 14980 19840 15008
rect 19484 14968 19490 14980
rect 19812 14952 19840 14980
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20732 15008 20760 15104
rect 24670 15036 24676 15088
rect 24728 15036 24734 15088
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20732 14980 20821 15008
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 21634 14968 21640 15020
rect 21692 15008 21698 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 21692 14980 22293 15008
rect 21692 14968 21698 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 22428 14980 23121 15008
rect 22428 14968 22434 14980
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 24486 14968 24492 15020
rect 24544 14968 24550 15020
rect 24688 15008 24716 15036
rect 24949 15011 25007 15017
rect 24949 15008 24961 15011
rect 24688 14980 24961 15008
rect 24949 14977 24961 14980
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 18187 14912 18460 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18690 14900 18696 14952
rect 18748 14940 18754 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 18748 14912 19349 14940
rect 18748 14900 18754 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 18049 14875 18107 14881
rect 18049 14841 18061 14875
rect 18095 14872 18107 14875
rect 18506 14872 18512 14884
rect 18095 14844 18512 14872
rect 18095 14841 18107 14844
rect 18049 14835 18107 14841
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 19352 14872 19380 14903
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 19610 14900 19616 14952
rect 19668 14900 19674 14952
rect 19794 14900 19800 14952
rect 19852 14900 19858 14952
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 22388 14912 22477 14940
rect 22388 14884 22416 14912
rect 22465 14909 22477 14912
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 23382 14900 23388 14952
rect 23440 14900 23446 14952
rect 19886 14872 19892 14884
rect 19352 14844 19892 14872
rect 19886 14832 19892 14844
rect 19944 14832 19950 14884
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 22094 14872 22100 14884
rect 22060 14844 22100 14872
rect 22060 14832 22066 14844
rect 22094 14832 22100 14844
rect 22152 14872 22158 14884
rect 22370 14872 22376 14884
rect 22152 14844 22376 14872
rect 22152 14832 22158 14844
rect 22370 14832 22376 14844
rect 22428 14832 22434 14884
rect 24578 14832 24584 14884
rect 24636 14872 24642 14884
rect 25225 14875 25283 14881
rect 25225 14872 25237 14875
rect 24636 14844 25237 14872
rect 24636 14832 24642 14844
rect 25225 14841 25237 14844
rect 25271 14841 25283 14875
rect 25225 14835 25283 14841
rect 18414 14804 18420 14816
rect 17972 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 20625 14807 20683 14813
rect 20625 14773 20637 14807
rect 20671 14804 20683 14807
rect 20714 14804 20720 14816
rect 20671 14776 20720 14804
rect 20671 14773 20683 14776
rect 20625 14767 20683 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21910 14764 21916 14816
rect 21968 14764 21974 14816
rect 25314 14764 25320 14816
rect 25372 14804 25378 14816
rect 25409 14807 25467 14813
rect 25409 14804 25421 14807
rect 25372 14776 25421 14804
rect 25372 14764 25378 14776
rect 25409 14773 25421 14776
rect 25455 14773 25467 14807
rect 25409 14767 25467 14773
rect 1104 14714 25852 14736
rect 1104 14662 4043 14714
rect 4095 14662 4107 14714
rect 4159 14662 4171 14714
rect 4223 14662 4235 14714
rect 4287 14662 4299 14714
rect 4351 14662 10230 14714
rect 10282 14662 10294 14714
rect 10346 14662 10358 14714
rect 10410 14662 10422 14714
rect 10474 14662 10486 14714
rect 10538 14662 16417 14714
rect 16469 14662 16481 14714
rect 16533 14662 16545 14714
rect 16597 14662 16609 14714
rect 16661 14662 16673 14714
rect 16725 14662 22604 14714
rect 22656 14662 22668 14714
rect 22720 14662 22732 14714
rect 22784 14662 22796 14714
rect 22848 14662 22860 14714
rect 22912 14662 25852 14714
rect 1104 14640 25852 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 2225 14603 2283 14609
rect 2225 14600 2237 14603
rect 1912 14572 2237 14600
rect 1912 14560 1918 14572
rect 2225 14569 2237 14572
rect 2271 14569 2283 14603
rect 2225 14563 2283 14569
rect 2406 14560 2412 14612
rect 2464 14560 2470 14612
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 3016 14572 3065 14600
rect 3016 14560 3022 14572
rect 3053 14569 3065 14572
rect 3099 14569 3111 14603
rect 11882 14600 11888 14612
rect 3053 14563 3111 14569
rect 5460 14572 11888 14600
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 2424 14405 2452 14560
rect 2866 14492 2872 14544
rect 2924 14492 2930 14544
rect 5350 14492 5356 14544
rect 5408 14492 5414 14544
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14365 2467 14399
rect 2409 14359 2467 14365
rect 2498 14356 2504 14408
rect 2556 14356 2562 14408
rect 2976 14396 3004 14427
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 5460 14464 5488 14572
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 13817 14603 13875 14609
rect 13817 14569 13829 14603
rect 13863 14600 13875 14603
rect 14274 14600 14280 14612
rect 13863 14572 14280 14600
rect 13863 14569 13875 14572
rect 13817 14563 13875 14569
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 18046 14600 18052 14612
rect 14660 14572 18052 14600
rect 9677 14535 9735 14541
rect 9677 14501 9689 14535
rect 9723 14532 9735 14535
rect 10042 14532 10048 14544
rect 9723 14504 10048 14532
rect 9723 14501 9735 14504
rect 9677 14495 9735 14501
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 14660 14532 14688 14572
rect 12406 14504 14688 14532
rect 3108 14436 5488 14464
rect 5813 14467 5871 14473
rect 3108 14424 3114 14436
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6362 14464 6368 14476
rect 5859 14436 6368 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 8202 14464 8208 14476
rect 8036 14436 8208 14464
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 2976 14368 3249 14396
rect 3237 14365 3249 14368
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 5534 14396 5540 14408
rect 3936 14368 5540 14396
rect 3936 14356 3942 14368
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 8036 14405 8064 14436
rect 8202 14424 8208 14436
rect 8260 14464 8266 14476
rect 12406 14464 12434 14504
rect 8260 14436 12434 14464
rect 14829 14467 14887 14473
rect 8260 14424 8266 14436
rect 14829 14433 14841 14467
rect 14875 14464 14887 14467
rect 15470 14464 15476 14476
rect 14875 14436 15476 14464
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 16666 14464 16672 14476
rect 16623 14436 16672 14464
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 4522 14328 4528 14340
rect 1596 14300 4528 14328
rect 1596 14269 1624 14300
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 4985 14331 5043 14337
rect 4985 14297 4997 14331
rect 5031 14328 5043 14331
rect 5074 14328 5080 14340
rect 5031 14300 5080 14328
rect 5031 14297 5043 14300
rect 4985 14291 5043 14297
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 5368 14300 6224 14328
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 5368 14260 5396 14300
rect 3292 14232 5396 14260
rect 5445 14263 5503 14269
rect 3292 14220 3298 14232
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5994 14260 6000 14272
rect 5491 14232 6000 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 6196 14260 6224 14300
rect 6362 14288 6368 14340
rect 6420 14288 6426 14340
rect 7834 14328 7840 14340
rect 7208 14300 7840 14328
rect 7208 14260 7236 14300
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 8168 14300 8309 14328
rect 8168 14288 8174 14300
rect 8297 14297 8309 14300
rect 8343 14297 8355 14331
rect 9876 14328 9904 14359
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 10560 14368 10609 14396
rect 10560 14356 10566 14368
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 16776 14405 16804 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 19978 14600 19984 14612
rect 18739 14572 19984 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 22465 14603 22523 14609
rect 21968 14572 22094 14600
rect 21968 14560 21974 14572
rect 18506 14492 18512 14544
rect 18564 14492 18570 14544
rect 20714 14424 20720 14476
rect 20772 14424 20778 14476
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14148 14368 14565 14396
rect 14148 14356 14154 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20438 14396 20444 14408
rect 19760 14368 20444 14396
rect 19760 14356 19766 14368
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 22066 14396 22094 14572
rect 22465 14569 22477 14603
rect 22511 14600 22523 14603
rect 23382 14600 23388 14612
rect 22511 14572 23388 14600
rect 22511 14569 22523 14572
rect 22465 14563 22523 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 23750 14560 23756 14612
rect 23808 14600 23814 14612
rect 24029 14603 24087 14609
rect 24029 14600 24041 14603
rect 23808 14572 24041 14600
rect 23808 14560 23814 14572
rect 24029 14569 24041 14572
rect 24075 14569 24087 14603
rect 24029 14563 24087 14569
rect 24486 14560 24492 14612
rect 24544 14600 24550 14612
rect 24949 14603 25007 14609
rect 24949 14600 24961 14603
rect 24544 14572 24961 14600
rect 24544 14560 24550 14572
rect 24949 14569 24961 14572
rect 24995 14569 25007 14603
rect 24949 14563 25007 14569
rect 25314 14560 25320 14612
rect 25372 14560 25378 14612
rect 25409 14603 25467 14609
rect 25409 14569 25421 14603
rect 25455 14600 25467 14603
rect 25455 14572 26004 14600
rect 25455 14569 25467 14572
rect 25409 14563 25467 14569
rect 23937 14535 23995 14541
rect 23937 14501 23949 14535
rect 23983 14532 23995 14535
rect 24578 14532 24584 14544
rect 23983 14504 24584 14532
rect 23983 14501 23995 14504
rect 23937 14495 23995 14501
rect 24578 14492 24584 14504
rect 24636 14532 24642 14544
rect 24673 14535 24731 14541
rect 24673 14532 24685 14535
rect 24636 14504 24685 14532
rect 24636 14492 24642 14504
rect 24673 14501 24685 14504
rect 24719 14532 24731 14535
rect 24762 14532 24768 14544
rect 24719 14504 24768 14532
rect 24719 14501 24731 14504
rect 24673 14495 24731 14501
rect 24762 14492 24768 14504
rect 24820 14492 24826 14544
rect 25332 14464 25360 14560
rect 25976 14544 26004 14572
rect 25958 14492 25964 14544
rect 26016 14492 26022 14544
rect 25148 14436 25360 14464
rect 22649 14399 22707 14405
rect 22649 14396 22661 14399
rect 22066 14368 22661 14396
rect 22649 14365 22661 14368
rect 22695 14365 22707 14399
rect 24489 14399 24547 14405
rect 24489 14396 24501 14399
rect 22649 14359 22707 14365
rect 23492 14368 24501 14396
rect 10318 14328 10324 14340
rect 9876 14300 10324 14328
rect 8297 14291 8355 14297
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 10873 14331 10931 14337
rect 10873 14328 10885 14331
rect 10836 14300 10885 14328
rect 10836 14288 10842 14300
rect 10873 14297 10885 14300
rect 10919 14297 10931 14331
rect 10873 14291 10931 14297
rect 11514 14288 11520 14340
rect 11572 14288 11578 14340
rect 13541 14331 13599 14337
rect 13541 14297 13553 14331
rect 13587 14328 13599 14331
rect 13630 14328 13636 14340
rect 13587 14300 13636 14328
rect 13587 14297 13599 14300
rect 13541 14291 13599 14297
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 15562 14288 15568 14340
rect 15620 14288 15626 14340
rect 18233 14331 18291 14337
rect 18233 14297 18245 14331
rect 18279 14328 18291 14331
rect 18414 14328 18420 14340
rect 18279 14300 18420 14328
rect 18279 14297 18291 14300
rect 18233 14291 18291 14297
rect 18414 14288 18420 14300
rect 18472 14288 18478 14340
rect 21358 14288 21364 14340
rect 21416 14288 21422 14340
rect 23492 14328 23520 14368
rect 24489 14365 24501 14368
rect 24535 14396 24547 14399
rect 24854 14396 24860 14408
rect 24535 14368 24860 14396
rect 24535 14365 24547 14368
rect 24489 14359 24547 14365
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 24946 14356 24952 14408
rect 25004 14356 25010 14408
rect 25148 14405 25176 14436
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14365 25191 14399
rect 25133 14359 25191 14365
rect 25225 14399 25283 14405
rect 25225 14365 25237 14399
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 22066 14300 23520 14328
rect 23569 14331 23627 14337
rect 6196 14232 7236 14260
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 11606 14260 11612 14272
rect 8628 14232 11612 14260
rect 8628 14220 8634 14232
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 15252 14232 16865 14260
rect 15252 14220 15258 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 22066 14260 22094 14300
rect 23569 14297 23581 14331
rect 23615 14328 23627 14331
rect 24670 14328 24676 14340
rect 23615 14300 24676 14328
rect 23615 14297 23627 14300
rect 23569 14291 23627 14297
rect 24670 14288 24676 14300
rect 24728 14288 24734 14340
rect 24964 14328 24992 14356
rect 25240 14328 25268 14359
rect 24964 14300 25268 14328
rect 20588 14232 22094 14260
rect 20588 14220 20594 14232
rect 22186 14220 22192 14272
rect 22244 14220 22250 14272
rect 1104 14170 25852 14192
rect 1104 14118 4703 14170
rect 4755 14118 4767 14170
rect 4819 14118 4831 14170
rect 4883 14118 4895 14170
rect 4947 14118 4959 14170
rect 5011 14118 10890 14170
rect 10942 14118 10954 14170
rect 11006 14118 11018 14170
rect 11070 14118 11082 14170
rect 11134 14118 11146 14170
rect 11198 14118 17077 14170
rect 17129 14118 17141 14170
rect 17193 14118 17205 14170
rect 17257 14118 17269 14170
rect 17321 14118 17333 14170
rect 17385 14118 23264 14170
rect 23316 14118 23328 14170
rect 23380 14118 23392 14170
rect 23444 14118 23456 14170
rect 23508 14118 23520 14170
rect 23572 14118 25852 14170
rect 1104 14096 25852 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 3050 14056 3056 14068
rect 1627 14028 3056 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14025 3203 14059
rect 3145 14019 3203 14025
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 3053 13923 3111 13929
rect 3053 13889 3065 13923
rect 3099 13920 3111 13923
rect 3160 13920 3188 14019
rect 3234 14016 3240 14068
rect 3292 14056 3298 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 3292 14028 3525 14056
rect 3292 14016 3298 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 3513 14019 3571 14025
rect 4614 14016 4620 14068
rect 4672 14016 4678 14068
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 7098 14056 7104 14068
rect 6656 14028 7104 14056
rect 3099 13892 3188 13920
rect 3605 13923 3663 13929
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4430 13920 4436 13932
rect 3651 13892 4436 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 4632 13920 4660 14016
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 6656 13988 6684 14028
rect 7098 14016 7104 14028
rect 7156 14056 7162 14068
rect 7156 14028 10180 14056
rect 7156 14016 7162 14028
rect 5592 13960 6684 13988
rect 5592 13948 5598 13960
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 4632 13892 5641 13920
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6656 13929 6684 13960
rect 7374 13948 7380 14000
rect 7432 13948 7438 14000
rect 8496 13929 8524 14028
rect 10042 13988 10048 14000
rect 9982 13960 10048 13988
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6052 13892 6561 13920
rect 6052 13880 6058 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 10152 13920 10180 14028
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10781 14059 10839 14065
rect 10781 14056 10793 14059
rect 10376 14028 10793 14056
rect 10376 14016 10382 14028
rect 10781 14025 10793 14028
rect 10827 14025 10839 14059
rect 10781 14019 10839 14025
rect 10873 14059 10931 14065
rect 10873 14025 10885 14059
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 10502 13948 10508 14000
rect 10560 13948 10566 14000
rect 10888 13988 10916 14019
rect 10796 13960 10916 13988
rect 10520 13920 10548 13948
rect 10796 13932 10824 13960
rect 10152 13892 10548 13920
rect 8481 13883 8539 13889
rect 10778 13880 10784 13932
rect 10836 13880 10842 13932
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11532 13920 11560 14019
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12342 14056 12348 14068
rect 12023 14028 12348 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 11992 13988 12020 14019
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12986 14056 12992 14068
rect 12584 14028 12992 14056
rect 12584 14016 12590 14028
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 15562 14016 15568 14068
rect 15620 14016 15626 14068
rect 15933 14059 15991 14065
rect 15933 14025 15945 14059
rect 15979 14056 15991 14059
rect 16298 14056 16304 14068
rect 15979 14028 16304 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 21542 14056 21548 14068
rect 21499 14028 21548 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 11848 13960 12020 13988
rect 14568 13960 16712 13988
rect 11848 13948 11854 13960
rect 11103 13892 11560 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 11606 13880 11612 13932
rect 11664 13920 11670 13932
rect 11664 13892 12434 13920
rect 11664 13880 11670 13892
rect 3786 13812 3792 13864
rect 3844 13812 3850 13864
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 5074 13852 5080 13864
rect 4939 13824 5080 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5350 13812 5356 13864
rect 5408 13812 5414 13864
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 10229 13855 10287 13861
rect 10229 13852 10241 13855
rect 9824 13824 10241 13852
rect 9824 13812 9830 13824
rect 10229 13821 10241 13824
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 11238 13852 11244 13864
rect 10367 13824 11244 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 11238 13812 11244 13824
rect 11296 13852 11302 13864
rect 11698 13852 11704 13864
rect 11296 13824 11704 13852
rect 11296 13812 11302 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 12406 13852 12434 13892
rect 12526 13880 12532 13932
rect 12584 13880 12590 13932
rect 14568 13929 14596 13960
rect 16684 13932 16712 13960
rect 20990 13948 20996 14000
rect 21048 13948 21054 14000
rect 24026 13948 24032 14000
rect 24084 13948 24090 14000
rect 24486 13948 24492 14000
rect 24544 13948 24550 14000
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14660 13852 14688 13883
rect 14734 13880 14740 13932
rect 14792 13880 14798 13932
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15286 13920 15292 13932
rect 14967 13892 15292 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15488 13892 15761 13920
rect 12406 13824 14688 13852
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 15488 13861 15516 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 16114 13880 16120 13932
rect 16172 13880 16178 13932
rect 16666 13880 16672 13932
rect 16724 13880 16730 13932
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13920 17739 13923
rect 17954 13920 17960 13932
rect 17727 13892 17960 13920
rect 17727 13889 17739 13892
rect 17681 13883 17739 13889
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14884 13824 15025 13852
rect 14884 13812 14890 13824
rect 15013 13821 15025 13824
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 19702 13812 19708 13864
rect 19760 13812 19766 13864
rect 19978 13812 19984 13864
rect 20036 13812 20042 13864
rect 23750 13812 23756 13864
rect 23808 13812 23814 13864
rect 25498 13812 25504 13864
rect 25556 13812 25562 13864
rect 5261 13787 5319 13793
rect 5261 13753 5273 13787
rect 5307 13784 5319 13787
rect 5368 13784 5396 13812
rect 6178 13784 6184 13796
rect 5307 13756 6184 13784
rect 5307 13753 5319 13756
rect 5261 13747 5319 13753
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 6546 13744 6552 13796
rect 6604 13744 6610 13796
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8168 13756 8524 13784
rect 8168 13744 8174 13756
rect 2866 13676 2872 13728
rect 2924 13676 2930 13728
rect 5350 13676 5356 13728
rect 5408 13676 5414 13728
rect 5442 13676 5448 13728
rect 5500 13676 5506 13728
rect 6564 13716 6592 13744
rect 8294 13716 8300 13728
rect 6564 13688 8300 13716
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8386 13676 8392 13728
rect 8444 13676 8450 13728
rect 8496 13716 8524 13756
rect 10686 13744 10692 13796
rect 10744 13784 10750 13796
rect 11606 13784 11612 13796
rect 10744 13756 11612 13784
rect 10744 13744 10750 13756
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 12250 13744 12256 13796
rect 12308 13784 12314 13796
rect 12308 13756 14872 13784
rect 12308 13744 12314 13756
rect 12158 13716 12164 13728
rect 8496 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12342 13676 12348 13728
rect 12400 13676 12406 13728
rect 14274 13676 14280 13728
rect 14332 13676 14338 13728
rect 14844 13716 14872 13756
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15289 13787 15347 13793
rect 15289 13784 15301 13787
rect 14976 13756 15301 13784
rect 14976 13744 14982 13756
rect 15289 13753 15301 13756
rect 15335 13753 15347 13787
rect 15289 13747 15347 13753
rect 16850 13744 16856 13796
rect 16908 13784 16914 13796
rect 17770 13784 17776 13796
rect 16908 13756 17776 13784
rect 16908 13744 16914 13756
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 19720 13784 19748 13812
rect 17880 13756 19748 13784
rect 17880 13728 17908 13756
rect 16758 13716 16764 13728
rect 14844 13688 16764 13716
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 17460 13688 17509 13716
rect 17460 13676 17466 13688
rect 17497 13685 17509 13688
rect 17543 13685 17555 13719
rect 17497 13679 17555 13685
rect 17862 13676 17868 13728
rect 17920 13676 17926 13728
rect 1104 13626 25852 13648
rect 1104 13574 4043 13626
rect 4095 13574 4107 13626
rect 4159 13574 4171 13626
rect 4223 13574 4235 13626
rect 4287 13574 4299 13626
rect 4351 13574 10230 13626
rect 10282 13574 10294 13626
rect 10346 13574 10358 13626
rect 10410 13574 10422 13626
rect 10474 13574 10486 13626
rect 10538 13574 16417 13626
rect 16469 13574 16481 13626
rect 16533 13574 16545 13626
rect 16597 13574 16609 13626
rect 16661 13574 16673 13626
rect 16725 13574 22604 13626
rect 22656 13574 22668 13626
rect 22720 13574 22732 13626
rect 22784 13574 22796 13626
rect 22848 13574 22860 13626
rect 22912 13574 25852 13626
rect 1104 13552 25852 13574
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 7374 13512 7380 13524
rect 6687 13484 7380 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 7490 13484 8708 13512
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 7190 13444 7196 13456
rect 6236 13416 7196 13444
rect 6236 13404 6242 13416
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 4338 13376 4344 13388
rect 3844 13348 4344 13376
rect 3844 13336 3850 13348
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 5902 13376 5908 13388
rect 5132 13348 5908 13376
rect 5132 13336 5138 13348
rect 5902 13336 5908 13348
rect 5960 13376 5966 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 5960 13348 6929 13376
rect 5960 13336 5966 13348
rect 6917 13345 6929 13348
rect 6963 13376 6975 13379
rect 7006 13376 7012 13388
rect 6963 13348 7012 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13308 3387 13311
rect 3375 13280 3832 13308
rect 3375 13277 3387 13280
rect 3329 13271 3387 13277
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13240 1547 13243
rect 3050 13240 3056 13252
rect 1535 13212 3056 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 3050 13200 3056 13212
rect 3108 13200 3114 13252
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 992 13144 1593 13172
rect 992 13132 998 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 3142 13132 3148 13184
rect 3200 13132 3206 13184
rect 3804 13181 3832 13280
rect 4522 13268 4528 13320
rect 4580 13268 4586 13320
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5350 13308 5356 13320
rect 4847 13280 5356 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7392 13308 7420 13339
rect 6871 13280 7420 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 4157 13243 4215 13249
rect 4157 13209 4169 13243
rect 4203 13240 4215 13243
rect 4540 13240 4568 13268
rect 4203 13212 5120 13240
rect 4203 13209 4215 13212
rect 4157 13203 4215 13209
rect 5092 13184 5120 13212
rect 7190 13200 7196 13252
rect 7248 13240 7254 13252
rect 7490 13240 7518 13484
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 8680 13444 8708 13484
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8812 13484 9045 13512
rect 8812 13472 8818 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 10594 13512 10600 13524
rect 9033 13475 9091 13481
rect 9876 13484 10600 13512
rect 9876 13444 9904 13484
rect 10594 13472 10600 13484
rect 10652 13472 10658 13524
rect 11149 13515 11207 13521
rect 11149 13481 11161 13515
rect 11195 13512 11207 13515
rect 12526 13512 12532 13524
rect 11195 13484 12532 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 12768 13484 13829 13512
rect 12768 13472 12774 13484
rect 13817 13481 13829 13484
rect 13863 13512 13875 13515
rect 16666 13512 16672 13524
rect 13863 13484 16672 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17678 13512 17684 13524
rect 16816 13484 17684 13512
rect 16816 13472 16822 13484
rect 17678 13472 17684 13484
rect 17736 13512 17742 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17736 13484 18153 13512
rect 17736 13472 17742 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 18598 13472 18604 13524
rect 18656 13472 18662 13524
rect 19889 13515 19947 13521
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 19978 13512 19984 13524
rect 19935 13484 19984 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20990 13472 20996 13524
rect 21048 13472 21054 13524
rect 21358 13472 21364 13524
rect 21416 13472 21422 13524
rect 24486 13472 24492 13524
rect 24544 13472 24550 13524
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 25133 13515 25191 13521
rect 25133 13512 25145 13515
rect 24912 13484 25145 13512
rect 24912 13472 24918 13484
rect 25133 13481 25145 13484
rect 25179 13481 25191 13515
rect 25133 13475 25191 13481
rect 8352 13416 8616 13444
rect 8680 13416 9904 13444
rect 8352 13404 8358 13416
rect 8110 13336 8116 13388
rect 8168 13336 8174 13388
rect 8588 13376 8616 13416
rect 8588 13348 9720 13376
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13308 8079 13311
rect 8386 13308 8392 13320
rect 8067 13280 8392 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9263 13280 9444 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 7248 13212 7518 13240
rect 7929 13243 7987 13249
rect 7248 13200 7254 13212
rect 7929 13209 7941 13243
rect 7975 13240 7987 13243
rect 7975 13212 8156 13240
rect 7975 13209 7987 13212
rect 7929 13203 7987 13209
rect 8128 13184 8156 13212
rect 3789 13175 3847 13181
rect 3789 13141 3801 13175
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 4522 13172 4528 13184
rect 4295 13144 4528 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 4614 13132 4620 13184
rect 4672 13132 4678 13184
rect 5074 13132 5080 13184
rect 5132 13132 5138 13184
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5350 13172 5356 13184
rect 5224 13144 5356 13172
rect 5224 13132 5230 13144
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 7558 13132 7564 13184
rect 7616 13132 7622 13184
rect 8110 13132 8116 13184
rect 8168 13132 8174 13184
rect 9416 13181 9444 13280
rect 9692 13240 9720 13348
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 9861 13379 9919 13385
rect 9861 13376 9873 13379
rect 9824 13348 9873 13376
rect 9824 13336 9830 13348
rect 9861 13345 9873 13348
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13376 10011 13379
rect 10042 13376 10048 13388
rect 9999 13348 10048 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10042 13336 10048 13348
rect 10100 13376 10106 13388
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 10100 13348 11805 13376
rect 10100 13336 10106 13348
rect 11793 13345 11805 13348
rect 11839 13376 11851 13379
rect 12434 13376 12440 13388
rect 11839 13348 12440 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12434 13336 12440 13348
rect 12492 13376 12498 13388
rect 13630 13376 13636 13388
rect 12492 13348 13636 13376
rect 12492 13336 12498 13348
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 14108 13348 16405 13376
rect 14108 13320 14136 13348
rect 16393 13345 16405 13348
rect 16439 13376 16451 13379
rect 17862 13376 17868 13388
rect 16439 13348 17868 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18616 13376 18644 13472
rect 20165 13447 20223 13453
rect 20165 13413 20177 13447
rect 20211 13413 20223 13447
rect 20165 13407 20223 13413
rect 18248 13348 18644 13376
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 12069 13311 12127 13317
rect 10836 13280 11744 13308
rect 10836 13268 10842 13280
rect 10686 13240 10692 13252
rect 9692 13212 10692 13240
rect 10686 13200 10692 13212
rect 10744 13240 10750 13252
rect 11517 13243 11575 13249
rect 11517 13240 11529 13243
rect 10744 13212 11529 13240
rect 10744 13200 10750 13212
rect 11517 13209 11529 13212
rect 11563 13209 11575 13243
rect 11716 13240 11744 13280
rect 12069 13277 12081 13311
rect 12115 13277 12127 13311
rect 12069 13271 12127 13277
rect 12084 13240 12112 13271
rect 13446 13268 13452 13320
rect 13504 13268 13510 13320
rect 14090 13268 14096 13320
rect 14148 13268 14154 13320
rect 16298 13268 16304 13320
rect 16356 13268 16362 13320
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 18248 13317 18276 13348
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 11716 13212 12112 13240
rect 11517 13203 11575 13209
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 12345 13243 12403 13249
rect 12345 13240 12357 13243
rect 12308 13212 12357 13240
rect 12308 13200 12314 13212
rect 12345 13209 12357 13212
rect 12391 13209 12403 13243
rect 12345 13203 12403 13209
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14369 13243 14427 13249
rect 14369 13240 14381 13243
rect 14332 13212 14381 13240
rect 14332 13200 14338 13212
rect 14369 13209 14381 13212
rect 14415 13209 14427 13243
rect 14369 13203 14427 13209
rect 15378 13200 15384 13252
rect 15436 13200 15442 13252
rect 16669 13243 16727 13249
rect 16669 13240 16681 13243
rect 16132 13212 16681 13240
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 9766 13132 9772 13184
rect 9824 13132 9830 13184
rect 11609 13175 11667 13181
rect 11609 13141 11621 13175
rect 11655 13172 11667 13175
rect 12434 13172 12440 13184
rect 11655 13144 12440 13172
rect 11655 13141 11667 13144
rect 11609 13135 11667 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 16132 13181 16160 13212
rect 16669 13209 16681 13212
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 17402 13200 17408 13252
rect 17460 13200 17466 13252
rect 18064 13240 18092 13268
rect 18616 13240 18644 13271
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20180 13308 20208 13407
rect 20254 13336 20260 13388
rect 20312 13376 20318 13388
rect 20622 13376 20628 13388
rect 20312 13348 20628 13376
rect 20312 13336 20318 13348
rect 20622 13336 20628 13348
rect 20680 13376 20686 13388
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 20680 13348 20729 13376
rect 20680 13336 20686 13348
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 20119 13280 20208 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 21174 13268 21180 13320
rect 21232 13268 21238 13320
rect 21542 13268 21548 13320
rect 21600 13268 21606 13320
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 24670 13268 24676 13320
rect 24728 13268 24734 13320
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13308 25283 13311
rect 25590 13308 25596 13320
rect 25271 13280 25596 13308
rect 25271 13277 25283 13280
rect 25225 13271 25283 13277
rect 18874 13240 18880 13252
rect 18064 13212 18880 13240
rect 18874 13200 18880 13212
rect 18932 13200 18938 13252
rect 20530 13200 20536 13252
rect 20588 13200 20594 13252
rect 24964 13240 24992 13271
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 25682 13268 25688 13320
rect 25740 13268 25746 13320
rect 25700 13240 25728 13268
rect 24964 13212 25728 13240
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13141 16175 13175
rect 16117 13135 16175 13141
rect 18414 13132 18420 13184
rect 18472 13132 18478 13184
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 18785 13175 18843 13181
rect 18785 13172 18797 13175
rect 18564 13144 18797 13172
rect 18564 13132 18570 13144
rect 18785 13141 18797 13144
rect 18831 13141 18843 13175
rect 18785 13135 18843 13141
rect 19245 13175 19303 13181
rect 19245 13141 19257 13175
rect 19291 13172 19303 13175
rect 19334 13172 19340 13184
rect 19291 13144 19340 13172
rect 19291 13141 19303 13144
rect 19245 13135 19303 13141
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 20625 13175 20683 13181
rect 20625 13141 20637 13175
rect 20671 13172 20683 13175
rect 21910 13172 21916 13184
rect 20671 13144 21916 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 23753 13175 23811 13181
rect 23753 13172 23765 13175
rect 23716 13144 23765 13172
rect 23716 13132 23722 13144
rect 23753 13141 23765 13144
rect 23799 13141 23811 13175
rect 23753 13135 23811 13141
rect 25406 13132 25412 13184
rect 25464 13132 25470 13184
rect 1104 13082 25852 13104
rect 1104 13030 4703 13082
rect 4755 13030 4767 13082
rect 4819 13030 4831 13082
rect 4883 13030 4895 13082
rect 4947 13030 4959 13082
rect 5011 13030 10890 13082
rect 10942 13030 10954 13082
rect 11006 13030 11018 13082
rect 11070 13030 11082 13082
rect 11134 13030 11146 13082
rect 11198 13030 17077 13082
rect 17129 13030 17141 13082
rect 17193 13030 17205 13082
rect 17257 13030 17269 13082
rect 17321 13030 17333 13082
rect 17385 13030 23264 13082
rect 23316 13030 23328 13082
rect 23380 13030 23392 13082
rect 23444 13030 23456 13082
rect 23508 13030 23520 13082
rect 23572 13030 25852 13082
rect 1104 13008 25852 13030
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 2924 12940 3096 12968
rect 2924 12928 2930 12940
rect 3068 12909 3096 12940
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 4525 12971 4583 12977
rect 4525 12968 4537 12971
rect 4488 12940 4537 12968
rect 4488 12928 4494 12940
rect 4525 12937 4537 12940
rect 4571 12968 4583 12971
rect 4706 12968 4712 12980
rect 4571 12940 4712 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6972 12940 7205 12968
rect 6972 12928 6978 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 7558 12928 7564 12980
rect 7616 12928 7622 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 8570 12968 8576 12980
rect 8527 12940 8576 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 10962 12968 10968 12980
rect 8720 12940 10968 12968
rect 8720 12928 8726 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 13262 12968 13268 12980
rect 11164 12940 13268 12968
rect 3053 12903 3111 12909
rect 3053 12869 3065 12903
rect 3099 12869 3111 12903
rect 4614 12900 4620 12912
rect 4278 12872 4620 12900
rect 3053 12863 3111 12869
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 7576 12900 7604 12928
rect 7392 12872 7604 12900
rect 2406 12792 2412 12844
rect 2464 12792 2470 12844
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 7392 12841 7420 12872
rect 7650 12860 7656 12912
rect 7708 12860 7714 12912
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 11164 12900 11192 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13446 12928 13452 12980
rect 13504 12928 13510 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 15013 12971 15071 12977
rect 13688 12940 14964 12968
rect 13688 12928 13694 12940
rect 8352 12872 11192 12900
rect 8352 12860 8358 12872
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 11296 12872 14013 12900
rect 11296 12860 11302 12872
rect 14001 12869 14013 12872
rect 14047 12900 14059 12903
rect 14553 12903 14611 12909
rect 14553 12900 14565 12903
rect 14047 12872 14565 12900
rect 14047 12869 14059 12872
rect 14001 12863 14059 12869
rect 14553 12869 14565 12872
rect 14599 12900 14611 12903
rect 14826 12900 14832 12912
rect 14599 12872 14832 12900
rect 14599 12869 14611 12872
rect 14553 12863 14611 12869
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 14936 12900 14964 12940
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 16114 12968 16120 12980
rect 15059 12940 16120 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 16298 12928 16304 12980
rect 16356 12968 16362 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16356 12940 16681 12968
rect 16356 12928 16362 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 17954 12928 17960 12980
rect 18012 12928 18018 12980
rect 20901 12971 20959 12977
rect 20901 12937 20913 12971
rect 20947 12968 20959 12971
rect 21174 12968 21180 12980
rect 20947 12940 21180 12968
rect 20947 12937 20959 12940
rect 20901 12931 20959 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21453 12971 21511 12977
rect 21453 12937 21465 12971
rect 21499 12968 21511 12971
rect 21542 12968 21548 12980
rect 21499 12940 21548 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 23106 12968 23112 12980
rect 22664 12940 23112 12968
rect 15194 12900 15200 12912
rect 14936 12872 15200 12900
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15565 12903 15623 12909
rect 15565 12900 15577 12903
rect 15344 12872 15577 12900
rect 15344 12860 15350 12872
rect 15565 12869 15577 12872
rect 15611 12900 15623 12903
rect 16022 12900 16028 12912
rect 15611 12872 16028 12900
rect 15611 12869 15623 12872
rect 15565 12863 15623 12869
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 16574 12860 16580 12912
rect 16632 12900 16638 12912
rect 17037 12903 17095 12909
rect 17037 12900 17049 12903
rect 16632 12872 17049 12900
rect 16632 12860 16638 12872
rect 17037 12869 17049 12872
rect 17083 12869 17095 12903
rect 17037 12863 17095 12869
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 18598 12900 18604 12912
rect 17543 12872 18604 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 19334 12860 19340 12912
rect 19392 12860 19398 12912
rect 20438 12860 20444 12912
rect 20496 12900 20502 12912
rect 22664 12900 22692 12940
rect 23106 12928 23112 12940
rect 23164 12968 23170 12980
rect 23750 12968 23756 12980
rect 23164 12940 23756 12968
rect 23164 12928 23170 12940
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 24394 12928 24400 12980
rect 24452 12928 24458 12980
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 24728 12940 25053 12968
rect 24728 12928 24734 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 20496 12872 22692 12900
rect 20496 12860 20502 12872
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7668 12832 7696 12860
rect 7607 12804 7696 12832
rect 7837 12835 7895 12841
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8110 12832 8116 12844
rect 7883 12804 8116 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10459 12804 10640 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 2884 12736 5028 12764
rect 2130 12656 2136 12708
rect 2188 12696 2194 12708
rect 2884 12696 2912 12736
rect 2188 12668 2912 12696
rect 2188 12656 2194 12668
rect 2225 12631 2283 12637
rect 2225 12597 2237 12631
rect 2271 12628 2283 12631
rect 2866 12628 2872 12640
rect 2271 12600 2872 12628
rect 2271 12597 2283 12600
rect 2225 12591 2283 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 4706 12588 4712 12640
rect 4764 12588 4770 12640
rect 5000 12628 5028 12736
rect 5074 12724 5080 12776
rect 5132 12764 5138 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 5132 12736 7665 12764
rect 5132 12724 5138 12736
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 9674 12764 9680 12776
rect 7653 12727 7711 12733
rect 7944 12736 9680 12764
rect 7944 12696 7972 12736
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9784 12764 9812 12792
rect 10502 12764 10508 12776
rect 9784 12736 10508 12764
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 9490 12696 9496 12708
rect 7484 12668 7972 12696
rect 8036 12668 9496 12696
rect 7484 12628 7512 12668
rect 5000 12600 7512 12628
rect 7834 12588 7840 12640
rect 7892 12588 7898 12640
rect 8036 12637 8064 12668
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 9692 12696 9720 12724
rect 10612 12696 10640 12804
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11422 12832 11428 12844
rect 11103 12804 11428 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12710 12832 12716 12844
rect 12483 12804 12716 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 13044 12804 13093 12832
rect 13044 12792 13050 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 11900 12764 11928 12792
rect 11440 12736 11928 12764
rect 11977 12767 12035 12773
rect 11440 12696 11468 12736
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12066 12764 12072 12776
rect 12023 12736 12072 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12342 12764 12348 12776
rect 12207 12736 12348 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 9692 12668 10640 12696
rect 10704 12668 11468 12696
rect 8021 12631 8079 12637
rect 8021 12597 8033 12631
rect 8067 12597 8079 12631
rect 8021 12591 8079 12597
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9858 12628 9864 12640
rect 9456 12600 9864 12628
rect 9456 12588 9462 12600
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10704 12637 10732 12668
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12989 12699 13047 12705
rect 12989 12696 13001 12699
rect 11940 12668 13001 12696
rect 11940 12656 11946 12668
rect 12989 12665 13001 12668
rect 13035 12665 13047 12699
rect 12989 12659 13047 12665
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12597 10747 12631
rect 10689 12591 10747 12597
rect 10870 12588 10876 12640
rect 10928 12588 10934 12640
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 11238 12628 11244 12640
rect 11020 12600 11244 12628
rect 11020 12588 11026 12600
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12628 11575 12631
rect 12434 12628 12440 12640
rect 11563 12600 12440 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 13096 12628 13124 12795
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 17402 12792 17408 12844
rect 17460 12792 17466 12844
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 18049 12835 18107 12841
rect 18049 12832 18061 12835
rect 17920 12804 18061 12832
rect 17920 12792 17926 12804
rect 18049 12801 18061 12804
rect 18095 12801 18107 12835
rect 20070 12832 20076 12844
rect 18049 12795 18107 12801
rect 19536 12804 20076 12832
rect 14458 12724 14464 12776
rect 14516 12724 14522 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15746 12764 15752 12776
rect 15252 12736 15752 12764
rect 15252 12724 15258 12736
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 17126 12724 17132 12776
rect 17184 12724 17190 12776
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12764 17371 12767
rect 17420 12764 17448 12792
rect 17359 12736 17448 12764
rect 17359 12733 17371 12736
rect 17313 12727 17371 12733
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19536 12764 19564 12804
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 20254 12792 20260 12844
rect 20312 12792 20318 12844
rect 22664 12841 22692 12872
rect 23658 12860 23664 12912
rect 23716 12860 23722 12912
rect 24578 12860 24584 12912
rect 24636 12860 24642 12912
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12832 25375 12835
rect 26050 12832 26056 12844
rect 25363 12804 26056 12832
rect 25363 12801 25375 12804
rect 25317 12795 25375 12801
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 18932 12736 19564 12764
rect 18932 12724 18938 12736
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20272 12764 20300 12792
rect 19852 12736 20300 12764
rect 19852 12724 19858 12736
rect 20346 12724 20352 12776
rect 20404 12764 20410 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20404 12736 20453 12764
rect 20404 12724 20410 12736
rect 20441 12733 20453 12736
rect 20487 12764 20499 12767
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20487 12736 21005 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20993 12733 21005 12736
rect 21039 12733 21051 12767
rect 20993 12727 21051 12733
rect 22922 12724 22928 12776
rect 22980 12724 22986 12776
rect 13262 12656 13268 12708
rect 13320 12696 13326 12708
rect 14277 12699 14335 12705
rect 14277 12696 14289 12699
rect 13320 12668 14289 12696
rect 13320 12656 13326 12668
rect 14277 12665 14289 12668
rect 14323 12696 14335 12699
rect 14829 12699 14887 12705
rect 14829 12696 14841 12699
rect 14323 12668 14841 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 14829 12665 14841 12668
rect 14875 12696 14887 12699
rect 14918 12696 14924 12708
rect 14875 12668 14924 12696
rect 14875 12665 14887 12668
rect 14829 12659 14887 12665
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 17773 12699 17831 12705
rect 17773 12665 17785 12699
rect 17819 12696 17831 12699
rect 18046 12696 18052 12708
rect 17819 12668 18052 12696
rect 17819 12665 17831 12668
rect 17773 12659 17831 12665
rect 17586 12628 17592 12640
rect 13096 12600 17592 12628
rect 17586 12588 17592 12600
rect 17644 12628 17650 12640
rect 17788 12628 17816 12659
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 20257 12699 20315 12705
rect 20257 12665 20269 12699
rect 20303 12696 20315 12699
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 20303 12668 20729 12696
rect 20303 12665 20315 12668
rect 20257 12659 20315 12665
rect 20717 12665 20729 12668
rect 20763 12696 20775 12699
rect 20806 12696 20812 12708
rect 20763 12668 20812 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 20806 12656 20812 12668
rect 20864 12696 20870 12708
rect 21269 12699 21327 12705
rect 21269 12696 21281 12699
rect 20864 12668 21281 12696
rect 20864 12656 20870 12668
rect 21269 12665 21281 12668
rect 21315 12665 21327 12699
rect 21269 12659 21327 12665
rect 24854 12656 24860 12708
rect 24912 12656 24918 12708
rect 25038 12656 25044 12708
rect 25096 12696 25102 12708
rect 25501 12699 25559 12705
rect 25501 12696 25513 12699
rect 25096 12668 25513 12696
rect 25096 12656 25102 12668
rect 25501 12665 25513 12668
rect 25547 12665 25559 12699
rect 25501 12659 25559 12665
rect 17644 12600 17816 12628
rect 17644 12588 17650 12600
rect 1104 12538 25852 12560
rect 1104 12486 4043 12538
rect 4095 12486 4107 12538
rect 4159 12486 4171 12538
rect 4223 12486 4235 12538
rect 4287 12486 4299 12538
rect 4351 12486 10230 12538
rect 10282 12486 10294 12538
rect 10346 12486 10358 12538
rect 10410 12486 10422 12538
rect 10474 12486 10486 12538
rect 10538 12486 16417 12538
rect 16469 12486 16481 12538
rect 16533 12486 16545 12538
rect 16597 12486 16609 12538
rect 16661 12486 16673 12538
rect 16725 12486 22604 12538
rect 22656 12486 22668 12538
rect 22720 12486 22732 12538
rect 22784 12486 22796 12538
rect 22848 12486 22860 12538
rect 22912 12486 25852 12538
rect 1104 12464 25852 12486
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 3108 12396 3157 12424
rect 3108 12384 3114 12396
rect 3145 12393 3157 12396
rect 3191 12424 3203 12427
rect 3234 12424 3240 12436
rect 3191 12396 3240 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 4890 12384 4896 12436
rect 4948 12424 4954 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 4948 12396 5733 12424
rect 4948 12384 4954 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 11514 12424 11520 12436
rect 5721 12387 5779 12393
rect 6380 12396 11520 12424
rect 2774 12316 2780 12368
rect 2832 12316 2838 12368
rect 2792 12288 2820 12316
rect 3878 12288 3884 12300
rect 2792 12260 3884 12288
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4706 12288 4712 12300
rect 4203 12260 4712 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 6380 12297 6408 12396
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12216 12396 12633 12424
rect 12216 12384 12222 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13630 12424 13636 12436
rect 13495 12396 13636 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 15378 12424 15384 12436
rect 14783 12396 15384 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 18233 12427 18291 12433
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 18322 12424 18328 12436
rect 18279 12396 18328 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19061 12427 19119 12433
rect 19061 12393 19073 12427
rect 19107 12424 19119 12427
rect 19426 12424 19432 12436
rect 19107 12396 19432 12424
rect 19107 12393 19119 12396
rect 19061 12387 19119 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 20346 12424 20352 12436
rect 19567 12396 20352 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 23845 12427 23903 12433
rect 23845 12393 23857 12427
rect 23891 12424 23903 12427
rect 23934 12424 23940 12436
rect 23891 12396 23940 12424
rect 23891 12393 23903 12396
rect 23845 12387 23903 12393
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 10870 12316 10876 12368
rect 10928 12316 10934 12368
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 12406 12328 12725 12356
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12257 6423 12291
rect 8570 12288 8576 12300
rect 6365 12251 6423 12257
rect 7484 12260 8576 12288
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 5534 12220 5540 12232
rect 5290 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 7484 12229 7512 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 10042 12288 10048 12300
rect 9456 12260 10048 12288
rect 9456 12248 9462 12260
rect 10042 12248 10048 12260
rect 10100 12288 10106 12300
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 10100 12260 10149 12288
rect 10100 12248 10106 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 10888 12288 10916 12316
rect 10744 12260 10916 12288
rect 11149 12291 11207 12297
rect 10744 12248 10750 12260
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 12406 12288 12434 12328
rect 12713 12325 12725 12328
rect 12759 12325 12771 12359
rect 12713 12319 12771 12325
rect 13262 12316 13268 12368
rect 13320 12316 13326 12368
rect 17037 12359 17095 12365
rect 17037 12325 17049 12359
rect 17083 12356 17095 12359
rect 17083 12328 18460 12356
rect 17083 12325 17095 12328
rect 17037 12319 17095 12325
rect 11195 12260 12434 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13044 12260 13676 12288
rect 13044 12248 13050 12260
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12121 1731 12155
rect 2958 12152 2964 12164
rect 2898 12124 2964 12152
rect 1673 12115 1731 12121
rect 1688 12084 1716 12115
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 7392 12152 7420 12183
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 7834 12220 7840 12232
rect 7791 12192 7840 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9732 12192 9965 12220
rect 9732 12180 9738 12192
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10836 12192 10885 12220
rect 10836 12180 10842 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 13648 12229 13676 12260
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17460 12260 17601 12288
rect 17460 12248 17466 12260
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 17678 12248 17684 12300
rect 17736 12248 17742 12300
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12492 12192 12909 12220
rect 12492 12180 12498 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 12897 12183 12955 12189
rect 13280 12192 13553 12220
rect 11054 12152 11060 12164
rect 3068 12124 3280 12152
rect 3068 12084 3096 12124
rect 1688 12056 3096 12084
rect 3252 12084 3280 12124
rect 5460 12124 7144 12152
rect 7392 12124 11060 12152
rect 5460 12084 5488 12124
rect 3252 12056 5488 12084
rect 5629 12087 5687 12093
rect 5629 12053 5641 12087
rect 5675 12084 5687 12087
rect 5810 12084 5816 12096
rect 5675 12056 5816 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 5810 12044 5816 12056
rect 5868 12084 5874 12096
rect 7116 12093 7144 12124
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 12158 12112 12164 12164
rect 12216 12112 12222 12164
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 13078 12152 13084 12164
rect 13035 12124 13084 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 5868 12056 6193 12084
rect 5868 12044 5874 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 7101 12087 7159 12093
rect 7101 12053 7113 12087
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 10042 12044 10048 12096
rect 10100 12044 10106 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 13280 12084 13308 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 14516 12192 14933 12220
rect 14516 12180 14522 12192
rect 14921 12189 14933 12192
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17696 12220 17724 12248
rect 18432 12229 18460 12328
rect 18874 12316 18880 12368
rect 18932 12316 18938 12368
rect 19306 12328 20668 12356
rect 18598 12248 18604 12300
rect 18656 12248 18662 12300
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 19306 12288 19334 12328
rect 18748 12260 19334 12288
rect 18748 12248 18754 12260
rect 20530 12248 20536 12300
rect 20588 12248 20594 12300
rect 20640 12288 20668 12328
rect 21910 12316 21916 12368
rect 21968 12356 21974 12368
rect 22281 12359 22339 12365
rect 22281 12356 22293 12359
rect 21968 12328 22293 12356
rect 21968 12316 21974 12328
rect 22281 12325 22293 12328
rect 22327 12325 22339 12359
rect 22281 12319 22339 12325
rect 23753 12359 23811 12365
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 24026 12356 24032 12368
rect 23799 12328 24032 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 24026 12316 24032 12328
rect 24084 12356 24090 12368
rect 24762 12356 24768 12368
rect 24084 12328 24768 12356
rect 24084 12316 24090 12328
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 23842 12288 23848 12300
rect 20640 12260 23848 12288
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24578 12248 24584 12300
rect 24636 12248 24642 12300
rect 17543 12192 17724 12220
rect 17865 12223 17923 12229
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 18616 12220 18644 12248
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 18616 12192 19441 12220
rect 17880 12152 17908 12183
rect 18616 12152 18644 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 20438 12180 20444 12232
rect 20496 12180 20502 12232
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 23658 12220 23664 12232
rect 23431 12192 23664 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 23658 12180 23664 12192
rect 23716 12220 23722 12232
rect 24596 12220 24624 12248
rect 23716 12192 24624 12220
rect 23716 12180 23722 12192
rect 20809 12155 20867 12161
rect 20809 12152 20821 12155
rect 17880 12124 18644 12152
rect 20272 12124 20821 12152
rect 11388 12056 13308 12084
rect 17405 12087 17463 12093
rect 11388 12044 11394 12056
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 17678 12084 17684 12096
rect 17451 12056 17684 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 20272 12093 20300 12124
rect 20809 12121 20821 12124
rect 20855 12121 20867 12155
rect 20809 12115 20867 12121
rect 21450 12112 21456 12164
rect 21508 12112 21514 12164
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 25958 12152 25964 12164
rect 22152 12124 25964 12152
rect 22152 12112 22158 12124
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 17920 12056 18061 12084
rect 17920 12044 17926 12056
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 20257 12087 20315 12093
rect 20257 12053 20269 12087
rect 20303 12053 20315 12087
rect 20257 12047 20315 12053
rect 1104 11994 25852 12016
rect 1104 11942 4703 11994
rect 4755 11942 4767 11994
rect 4819 11942 4831 11994
rect 4883 11942 4895 11994
rect 4947 11942 4959 11994
rect 5011 11942 10890 11994
rect 10942 11942 10954 11994
rect 11006 11942 11018 11994
rect 11070 11942 11082 11994
rect 11134 11942 11146 11994
rect 11198 11942 17077 11994
rect 17129 11942 17141 11994
rect 17193 11942 17205 11994
rect 17257 11942 17269 11994
rect 17321 11942 17333 11994
rect 17385 11942 23264 11994
rect 23316 11942 23328 11994
rect 23380 11942 23392 11994
rect 23444 11942 23456 11994
rect 23508 11942 23520 11994
rect 23572 11942 25852 11994
rect 1104 11920 25852 11942
rect 2406 11840 2412 11892
rect 2464 11840 2470 11892
rect 4522 11840 4528 11892
rect 4580 11840 4586 11892
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 3050 11772 3056 11824
rect 3108 11772 3114 11824
rect 4632 11812 4660 11843
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 6178 11880 6184 11892
rect 5132 11852 6184 11880
rect 5132 11840 5138 11852
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7558 11880 7564 11892
rect 7515 11852 7564 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 8846 11880 8852 11892
rect 8435 11852 8852 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 8404 11812 8432 11843
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 11330 11840 11336 11892
rect 11388 11840 11394 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11698 11880 11704 11892
rect 11572 11852 11704 11880
rect 11572 11840 11578 11852
rect 11698 11840 11704 11852
rect 11756 11880 11762 11892
rect 11756 11852 18368 11880
rect 11756 11840 11762 11852
rect 4278 11784 4660 11812
rect 4724 11784 7420 11812
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1854 11636 1860 11688
rect 1912 11676 1918 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1912 11648 1961 11676
rect 1912 11636 1918 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 2774 11676 2780 11688
rect 1949 11639 2007 11645
rect 2240 11648 2780 11676
rect 1394 11568 1400 11620
rect 1452 11608 1458 11620
rect 2240 11608 2268 11648
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 4724 11676 4752 11784
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 4847 11716 5396 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5368 11685 5396 11716
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6880 11716 7297 11744
rect 6880 11704 6886 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 2884 11648 4752 11676
rect 4893 11679 4951 11685
rect 1452 11580 2268 11608
rect 1452 11568 1458 11580
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 2884 11608 2912 11648
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 5353 11679 5411 11685
rect 4939 11648 5304 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 2372 11580 2912 11608
rect 2372 11568 2378 11580
rect 5074 11568 5080 11620
rect 5132 11608 5138 11620
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 5132 11580 5181 11608
rect 5132 11568 5138 11580
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5276 11608 5304 11648
rect 5353 11645 5365 11679
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 5920 11608 5948 11704
rect 7392 11676 7420 11784
rect 7484 11784 8432 11812
rect 7484 11753 7512 11784
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7800 11716 8125 11744
rect 7800 11704 7806 11716
rect 8113 11713 8125 11716
rect 8159 11744 8171 11747
rect 8202 11744 8208 11756
rect 8159 11716 8208 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9600 11753 9628 11840
rect 18340 11824 18368 11852
rect 20438 11840 20444 11892
rect 20496 11840 20502 11892
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 21821 11883 21879 11889
rect 21821 11849 21833 11883
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 9674 11772 9680 11824
rect 9732 11812 9738 11824
rect 10873 11815 10931 11821
rect 10873 11812 10885 11815
rect 9732 11784 10885 11812
rect 9732 11772 9738 11784
rect 10873 11781 10885 11784
rect 10919 11781 10931 11815
rect 10873 11775 10931 11781
rect 10980 11784 12388 11812
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 8294 11676 8300 11688
rect 7392 11648 8300 11676
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 6270 11608 6276 11620
rect 5276 11580 6276 11608
rect 5169 11571 5227 11577
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 10980 11608 11008 11784
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11514 11704 11520 11756
rect 11572 11704 11578 11756
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12066 11744 12072 11756
rect 11940 11716 12072 11744
rect 11940 11704 11946 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11977 11679 12035 11685
rect 11103 11648 11192 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 6564 11580 11008 11608
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 6564 11540 6592 11580
rect 1627 11512 6592 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 6638 11500 6644 11552
rect 6696 11500 6702 11552
rect 9398 11500 9404 11552
rect 9456 11500 9462 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10744 11512 10885 11540
rect 10744 11500 10750 11512
rect 10873 11509 10885 11512
rect 10919 11509 10931 11543
rect 11164 11540 11192 11648
rect 11977 11645 11989 11679
rect 12023 11676 12035 11679
rect 12268 11676 12296 11707
rect 12023 11648 12296 11676
rect 12360 11676 12388 11784
rect 18322 11772 18328 11824
rect 18380 11772 18386 11824
rect 20346 11772 20352 11824
rect 20404 11772 20410 11824
rect 20456 11812 20484 11840
rect 21836 11812 21864 11843
rect 22370 11840 22376 11892
rect 22428 11880 22434 11892
rect 23750 11880 23756 11892
rect 22428 11852 23756 11880
rect 22428 11840 22434 11852
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 24857 11883 24915 11889
rect 24857 11849 24869 11883
rect 24903 11880 24915 11883
rect 25130 11880 25136 11892
rect 24903 11852 25136 11880
rect 24903 11849 24915 11852
rect 24857 11843 24915 11849
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 25314 11840 25320 11892
rect 25372 11840 25378 11892
rect 20456 11784 21864 11812
rect 22189 11815 22247 11821
rect 22189 11781 22201 11815
rect 22235 11812 22247 11815
rect 25332 11812 25360 11840
rect 22235 11784 25360 11812
rect 22235 11781 22247 11784
rect 22189 11775 22247 11781
rect 15378 11704 15384 11756
rect 15436 11704 15442 11756
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17586 11744 17592 11756
rect 17359 11716 17592 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17586 11704 17592 11716
rect 17644 11704 17650 11756
rect 20364 11744 20392 11772
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 20364 11716 20913 11744
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 21637 11747 21695 11753
rect 21637 11713 21649 11747
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 21361 11679 21419 11685
rect 12360 11648 18828 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 18800 11620 18828 11648
rect 21361 11645 21373 11679
rect 21407 11676 21419 11679
rect 21652 11676 21680 11707
rect 24762 11704 24768 11756
rect 24820 11704 24826 11756
rect 21407 11648 21680 11676
rect 21407 11645 21419 11648
rect 21361 11639 21419 11645
rect 22278 11636 22284 11688
rect 22336 11636 22342 11688
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 11793 11611 11851 11617
rect 11793 11608 11805 11611
rect 11664 11580 11805 11608
rect 11664 11568 11670 11580
rect 11793 11577 11805 11580
rect 11839 11577 11851 11611
rect 11793 11571 11851 11577
rect 12069 11611 12127 11617
rect 12069 11577 12081 11611
rect 12115 11608 12127 11611
rect 12158 11608 12164 11620
rect 12115 11580 12164 11608
rect 12115 11577 12127 11580
rect 12069 11571 12127 11577
rect 11514 11540 11520 11552
rect 11164 11512 11520 11540
rect 10873 11503 10931 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11808 11540 11836 11571
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 18506 11608 18512 11620
rect 12406 11580 18512 11608
rect 12406 11540 12434 11580
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 18782 11568 18788 11620
rect 18840 11568 18846 11620
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 20864 11580 21189 11608
rect 20864 11568 20870 11580
rect 21177 11577 21189 11580
rect 21223 11577 21235 11611
rect 21177 11571 21235 11577
rect 11808 11512 12434 11540
rect 15473 11543 15531 11549
rect 15473 11509 15485 11543
rect 15519 11540 15531 11543
rect 15838 11540 15844 11552
rect 15519 11512 15844 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 17497 11543 17555 11549
rect 17497 11509 17509 11543
rect 17543 11540 17555 11543
rect 17954 11540 17960 11552
rect 17543 11512 17960 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 17954 11500 17960 11512
rect 18012 11500 18018 11552
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 22388 11540 22416 11639
rect 23750 11636 23756 11688
rect 23808 11676 23814 11688
rect 24949 11679 25007 11685
rect 24949 11676 24961 11679
rect 23808 11648 24961 11676
rect 23808 11636 23814 11648
rect 24949 11645 24961 11648
rect 24995 11645 25007 11679
rect 24949 11639 25007 11645
rect 21416 11512 22416 11540
rect 21416 11500 21422 11512
rect 24394 11500 24400 11552
rect 24452 11500 24458 11552
rect 1104 11450 25852 11472
rect 1104 11398 4043 11450
rect 4095 11398 4107 11450
rect 4159 11398 4171 11450
rect 4223 11398 4235 11450
rect 4287 11398 4299 11450
rect 4351 11398 10230 11450
rect 10282 11398 10294 11450
rect 10346 11398 10358 11450
rect 10410 11398 10422 11450
rect 10474 11398 10486 11450
rect 10538 11398 16417 11450
rect 16469 11398 16481 11450
rect 16533 11398 16545 11450
rect 16597 11398 16609 11450
rect 16661 11398 16673 11450
rect 16725 11398 22604 11450
rect 22656 11398 22668 11450
rect 22720 11398 22732 11450
rect 22784 11398 22796 11450
rect 22848 11398 22860 11450
rect 22912 11398 25852 11450
rect 1104 11376 25852 11398
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 3252 11308 4445 11336
rect 3252 11212 3280 11308
rect 4433 11305 4445 11308
rect 4479 11305 4491 11339
rect 4433 11299 4491 11305
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3234 11200 3240 11212
rect 3099 11172 3240 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 4448 11200 4476 11299
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4580 11308 4997 11336
rect 4580 11296 4586 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 6546 11296 6552 11348
rect 6604 11296 6610 11348
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 6822 11336 6828 11348
rect 6779 11308 6828 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 9398 11345 9404 11348
rect 9388 11339 9404 11345
rect 7248 11308 8708 11336
rect 7248 11296 7254 11308
rect 6564 11268 6592 11296
rect 7377 11271 7435 11277
rect 7377 11268 7389 11271
rect 6564 11240 7389 11268
rect 7377 11237 7389 11240
rect 7423 11237 7435 11271
rect 7377 11231 7435 11237
rect 8294 11228 8300 11280
rect 8352 11228 8358 11280
rect 5718 11200 5724 11212
rect 4448 11172 4936 11200
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 4522 11132 4528 11144
rect 4387 11104 4528 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 4908 11141 4936 11172
rect 5644 11172 5724 11200
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5442 11092 5448 11144
rect 5500 11092 5506 11144
rect 5644 11141 5672 11172
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 8680 11200 8708 11308
rect 9388 11305 9400 11339
rect 9388 11299 9404 11305
rect 9398 11296 9404 11299
rect 9456 11296 9462 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10100 11308 10885 11336
rect 10100 11296 10106 11308
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 13722 11336 13728 11348
rect 10919 11308 13728 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14240 11308 14565 11336
rect 14240 11296 14246 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 12618 11268 12624 11280
rect 11256 11240 12624 11268
rect 11256 11200 11284 11240
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 13906 11268 13912 11280
rect 13136 11240 13912 11268
rect 13136 11228 13142 11240
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 14568 11268 14596 11299
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14792 11308 15485 11336
rect 14792 11296 14798 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 17773 11339 17831 11345
rect 17773 11305 17785 11339
rect 17819 11336 17831 11339
rect 18874 11336 18880 11348
rect 17819 11308 18880 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 22833 11339 22891 11345
rect 22833 11305 22845 11339
rect 22879 11336 22891 11339
rect 22922 11336 22928 11348
rect 22879 11308 22928 11336
rect 22879 11305 22891 11308
rect 22833 11299 22891 11305
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 24394 11296 24400 11348
rect 24452 11296 24458 11348
rect 24762 11296 24768 11348
rect 24820 11336 24826 11348
rect 25317 11339 25375 11345
rect 25317 11336 25329 11339
rect 24820 11308 25329 11336
rect 24820 11296 24826 11308
rect 25317 11305 25329 11308
rect 25363 11305 25375 11339
rect 25317 11299 25375 11305
rect 15289 11271 15347 11277
rect 15289 11268 15301 11271
rect 14568 11240 15301 11268
rect 15289 11237 15301 11240
rect 15335 11237 15347 11271
rect 17681 11271 17739 11277
rect 15289 11231 15347 11237
rect 15768 11240 16344 11268
rect 6604 11172 7696 11200
rect 8680 11172 11284 11200
rect 6604 11160 6610 11172
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 6457 11135 6515 11141
rect 5675 11104 6408 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 2130 11064 2136 11076
rect 1535 11036 2136 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 4154 11064 4160 11076
rect 3651 11036 4160 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 6380 11064 6408 11104
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6638 11132 6644 11144
rect 6503 11104 6644 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7282 11132 7288 11144
rect 6972 11104 7288 11132
rect 6972 11092 6978 11104
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7558 11064 7564 11076
rect 6380 11036 7564 11064
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 7668 11064 7696 11172
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11606 11200 11612 11212
rect 11388 11172 11612 11200
rect 11388 11160 11394 11172
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 13354 11200 13360 11212
rect 12406 11172 13360 11200
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8662 11132 8668 11144
rect 7975 11104 8668 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8812 11104 9137 11132
rect 8812 11092 8818 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 11054 11132 11060 11144
rect 10534 11104 11060 11132
rect 9125 11095 9183 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 12406 11064 12434 11172
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14476 11172 15025 11200
rect 14476 11141 14504 11172
rect 15013 11169 15025 11172
rect 15059 11200 15071 11203
rect 15768 11200 15796 11240
rect 15059 11172 15796 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15838 11160 15844 11212
rect 15896 11200 15902 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15896 11172 16037 11200
rect 15896 11160 15902 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16206 11200 16212 11212
rect 16163 11172 16212 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15746 11132 15752 11144
rect 14608 11104 15752 11132
rect 14608 11092 14614 11104
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 16316 11141 16344 11240
rect 17681 11237 17693 11271
rect 17727 11268 17739 11271
rect 17954 11268 17960 11280
rect 17727 11240 17960 11268
rect 17727 11237 17739 11240
rect 17681 11231 17739 11237
rect 17954 11228 17960 11240
rect 18012 11268 18018 11280
rect 18141 11271 18199 11277
rect 18141 11268 18153 11271
rect 18012 11240 18153 11268
rect 18012 11228 18018 11240
rect 18141 11237 18153 11240
rect 18187 11237 18199 11271
rect 18141 11231 18199 11237
rect 20257 11271 20315 11277
rect 20257 11237 20269 11271
rect 20303 11268 20315 11271
rect 20303 11240 21312 11268
rect 20303 11237 20315 11240
rect 20257 11231 20315 11237
rect 17862 11200 17868 11212
rect 17420 11172 17868 11200
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16347 11104 16896 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 7668 11036 9812 11064
rect 1578 10956 1584 11008
rect 1636 10956 1642 11008
rect 4801 10999 4859 11005
rect 4801 10965 4813 10999
rect 4847 10996 4859 10999
rect 5074 10996 5080 11008
rect 4847 10968 5080 10996
rect 4847 10965 4859 10968
rect 4801 10959 4859 10965
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5350 10956 5356 11008
rect 5408 10956 5414 11008
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 8386 10956 8392 11008
rect 8444 10956 8450 11008
rect 9784 10996 9812 11036
rect 10704 11036 12434 11064
rect 15948 11064 15976 11095
rect 16758 11064 16764 11076
rect 15948 11036 16764 11064
rect 10704 10996 10732 11036
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 9784 10968 10732 10996
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 12434 10996 12440 11008
rect 11204 10968 12440 10996
rect 11204 10956 11210 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14734 10996 14740 11008
rect 14332 10968 14740 10996
rect 14332 10956 14338 10968
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 16482 10956 16488 11008
rect 16540 10956 16546 11008
rect 16868 10996 16896 11104
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17420 11064 17448 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 18371 11172 18644 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 18616 11141 18644 11172
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20588 11172 20821 11200
rect 20588 11160 20594 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 18840 11104 20637 11132
rect 18840 11092 18846 11104
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 20824 11132 20852 11163
rect 21174 11132 21180 11144
rect 20824 11104 21180 11132
rect 20625 11095 20683 11101
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 21284 11141 21312 11240
rect 24026 11228 24032 11280
rect 24084 11228 24090 11280
rect 23658 11160 23664 11212
rect 23716 11160 23722 11212
rect 24121 11203 24179 11209
rect 24121 11169 24133 11203
rect 24167 11169 24179 11203
rect 24121 11163 24179 11169
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 23014 11092 23020 11144
rect 23072 11092 23078 11144
rect 18708 11064 18736 11092
rect 17368 11036 17448 11064
rect 17972 11036 18736 11064
rect 20717 11067 20775 11073
rect 17368 11024 17374 11036
rect 17972 10996 18000 11036
rect 20717 11033 20729 11067
rect 20763 11064 20775 11067
rect 21910 11064 21916 11076
rect 20763 11036 21916 11064
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 21910 11024 21916 11036
rect 21968 11064 21974 11076
rect 22094 11064 22100 11076
rect 21968 11036 22100 11064
rect 21968 11024 21974 11036
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 24136 11064 24164 11163
rect 24412 11132 24440 11296
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24412 11104 24593 11132
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25501 11135 25559 11141
rect 25501 11101 25513 11135
rect 25547 11132 25559 11135
rect 25547 11104 26004 11132
rect 25547 11101 25559 11104
rect 25501 11095 25559 11101
rect 24872 11064 24900 11095
rect 25976 11076 26004 11104
rect 24136 11036 24900 11064
rect 25958 11024 25964 11076
rect 26016 11024 26022 11076
rect 16868 10968 18000 10996
rect 18414 10956 18420 11008
rect 18472 10956 18478 11008
rect 21082 10956 21088 11008
rect 21140 10956 21146 11008
rect 24394 10956 24400 11008
rect 24452 10956 24458 11008
rect 24670 10956 24676 11008
rect 24728 10956 24734 11008
rect 1104 10906 25852 10928
rect 1104 10854 4703 10906
rect 4755 10854 4767 10906
rect 4819 10854 4831 10906
rect 4883 10854 4895 10906
rect 4947 10854 4959 10906
rect 5011 10854 10890 10906
rect 10942 10854 10954 10906
rect 11006 10854 11018 10906
rect 11070 10854 11082 10906
rect 11134 10854 11146 10906
rect 11198 10854 17077 10906
rect 17129 10854 17141 10906
rect 17193 10854 17205 10906
rect 17257 10854 17269 10906
rect 17321 10854 17333 10906
rect 17385 10854 23264 10906
rect 23316 10854 23328 10906
rect 23380 10854 23392 10906
rect 23444 10854 23456 10906
rect 23508 10854 23520 10906
rect 23572 10854 25852 10906
rect 1104 10832 25852 10854
rect 8754 10792 8760 10804
rect 7668 10764 8760 10792
rect 5534 10724 5540 10736
rect 4724 10696 5540 10724
rect 1486 10616 1492 10668
rect 1544 10616 1550 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1912 10560 1961 10588
rect 1912 10548 1918 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2700 10588 2728 10619
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4724 10665 4752 10696
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 5997 10727 6055 10733
rect 5997 10724 6009 10727
rect 5960 10696 6009 10724
rect 5960 10684 5966 10696
rect 5997 10693 6009 10696
rect 6043 10693 6055 10727
rect 5997 10687 6055 10693
rect 6638 10684 6644 10736
rect 6696 10684 6702 10736
rect 7190 10684 7196 10736
rect 7248 10684 7254 10736
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4212 10628 4537 10656
rect 4212 10616 4218 10628
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 2455 10560 2728 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2314 10480 2320 10532
rect 2372 10480 2378 10532
rect 4632 10520 4660 10619
rect 4890 10616 4896 10668
rect 4948 10616 4954 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5074 10656 5080 10668
rect 5031 10628 5080 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 5000 10588 5028 10619
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5350 10616 5356 10668
rect 5408 10616 5414 10668
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 6656 10656 6684 10684
rect 5776 10628 6684 10656
rect 6733 10659 6791 10665
rect 5776 10616 5782 10628
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7208 10656 7236 10684
rect 6779 10628 7236 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 4856 10560 5028 10588
rect 5445 10591 5503 10597
rect 4856 10548 4862 10560
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 5491 10560 6009 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5997 10557 6009 10560
rect 6043 10588 6055 10591
rect 6043 10560 6776 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6748 10532 6776 10560
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7668 10597 7696 10764
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9674 10792 9680 10804
rect 9447 10764 9680 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 10134 10792 10140 10804
rect 9732 10764 10140 10792
rect 9732 10752 9738 10764
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10836 10764 10885 10792
rect 10836 10752 10842 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 11882 10752 11888 10804
rect 11940 10792 11946 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 11940 10764 12633 10792
rect 11940 10752 11946 10764
rect 12621 10761 12633 10764
rect 12667 10792 12679 10795
rect 18046 10792 18052 10804
rect 12667 10764 12940 10792
rect 12667 10761 12679 10764
rect 12621 10755 12679 10761
rect 8478 10684 8484 10736
rect 8536 10684 8542 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12912 10733 12940 10764
rect 13556 10764 18052 10792
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 12124 10696 12725 10724
rect 12124 10684 12130 10696
rect 12713 10693 12725 10696
rect 12759 10693 12771 10727
rect 12713 10687 12771 10693
rect 12897 10727 12955 10733
rect 12897 10693 12909 10727
rect 12943 10693 12955 10727
rect 12897 10687 12955 10693
rect 13556 10668 13584 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 18601 10795 18659 10801
rect 18601 10761 18613 10795
rect 18647 10792 18659 10795
rect 18690 10792 18696 10804
rect 18647 10764 18696 10792
rect 18647 10761 18659 10764
rect 18601 10755 18659 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 18785 10795 18843 10801
rect 18785 10761 18797 10795
rect 18831 10761 18843 10795
rect 18785 10755 18843 10761
rect 13998 10684 14004 10736
rect 14056 10724 14062 10736
rect 17218 10724 17224 10736
rect 14056 10696 15976 10724
rect 14056 10684 14062 10696
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9548 10628 9597 10656
rect 9548 10616 9554 10628
rect 9585 10625 9597 10628
rect 9631 10656 9643 10659
rect 13538 10656 13544 10668
rect 9631 10628 13544 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7156 10560 7665 10588
rect 7156 10548 7162 10560
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 7926 10548 7932 10600
rect 7984 10548 7990 10600
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 12032 10560 12173 10588
rect 12032 10548 12038 10560
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 13648 10588 13676 10619
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 14461 10660 14519 10665
rect 14384 10659 14519 10660
rect 14384 10656 14473 10659
rect 13780 10632 14473 10656
rect 13780 10628 14412 10632
rect 13780 10616 13786 10628
rect 14461 10625 14473 10632
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 15838 10616 15844 10668
rect 15896 10616 15902 10668
rect 15948 10665 15976 10696
rect 16868 10696 17224 10724
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16022 10616 16028 10668
rect 16080 10616 16086 10668
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16868 10665 16896 10696
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 18800 10724 18828 10755
rect 18874 10752 18880 10804
rect 18932 10752 18938 10804
rect 21082 10792 21088 10804
rect 20088 10764 21088 10792
rect 18354 10696 18828 10724
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 16172 10628 16221 10656
rect 16172 10616 16178 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 18892 10656 18920 10752
rect 20088 10733 20116 10764
rect 21082 10752 21088 10764
rect 21140 10752 21146 10804
rect 21821 10795 21879 10801
rect 21821 10761 21833 10795
rect 21867 10761 21879 10795
rect 24394 10792 24400 10804
rect 21821 10755 21879 10761
rect 23584 10764 24400 10792
rect 20073 10727 20131 10733
rect 20073 10693 20085 10727
rect 20119 10693 20131 10727
rect 21836 10724 21864 10755
rect 23584 10733 23612 10764
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 21298 10696 21864 10724
rect 23569 10727 23627 10733
rect 20073 10687 20131 10693
rect 23569 10693 23581 10727
rect 23615 10693 23627 10727
rect 23569 10687 23627 10693
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18892 10628 18981 10656
rect 16853 10619 16911 10625
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 23106 10616 23112 10668
rect 23164 10656 23170 10668
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 23164 10628 23305 10656
rect 23164 10616 23170 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 24670 10616 24676 10668
rect 24728 10616 24734 10668
rect 25225 10659 25283 10665
rect 25225 10625 25237 10659
rect 25271 10656 25283 10659
rect 25774 10656 25780 10668
rect 25271 10628 25780 10656
rect 25271 10625 25283 10628
rect 25225 10619 25283 10625
rect 25774 10616 25780 10628
rect 25832 10616 25838 10668
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 13648 10560 14749 10588
rect 12161 10551 12219 10557
rect 14737 10557 14749 10560
rect 14783 10588 14795 10591
rect 14783 10560 15056 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 5813 10523 5871 10529
rect 4632 10492 5764 10520
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 992 10424 1593 10452
rect 992 10412 998 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2464 10424 2513 10452
rect 2464 10412 2470 10424
rect 2501 10421 2513 10424
rect 2547 10421 2559 10455
rect 2501 10415 2559 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 3568 10424 4261 10452
rect 3568 10412 3574 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 5736 10452 5764 10492
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 6086 10520 6092 10532
rect 5859 10492 6092 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 6086 10480 6092 10492
rect 6144 10520 6150 10532
rect 6546 10520 6552 10532
rect 6144 10492 6552 10520
rect 6144 10480 6150 10492
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 6788 10492 7205 10520
rect 6788 10480 6794 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7193 10483 7251 10489
rect 11606 10480 11612 10532
rect 11664 10520 11670 10532
rect 12526 10520 12532 10532
rect 11664 10492 12532 10520
rect 11664 10480 11670 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 6822 10452 6828 10464
rect 5736 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6914 10412 6920 10464
rect 6972 10412 6978 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 12894 10452 12900 10464
rect 7800 10424 12900 10452
rect 7800 10412 7806 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13078 10412 13084 10464
rect 13136 10412 13142 10464
rect 13722 10412 13728 10464
rect 13780 10412 13786 10464
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10452 14151 10455
rect 14550 10452 14556 10464
rect 14139 10424 14556 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 15028 10452 15056 10560
rect 15286 10548 15292 10600
rect 15344 10548 15350 10600
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10588 15623 10591
rect 17129 10591 17187 10597
rect 17129 10588 17141 10591
rect 15611 10560 17141 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 17129 10557 17141 10560
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 19794 10588 19800 10600
rect 17276 10560 19800 10588
rect 17276 10548 17282 10560
rect 19794 10548 19800 10560
rect 19852 10548 19858 10600
rect 22741 10591 22799 10597
rect 22741 10557 22753 10591
rect 22787 10588 22799 10591
rect 23658 10588 23664 10600
rect 22787 10560 23664 10588
rect 22787 10557 22799 10560
rect 22741 10551 22799 10557
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 16298 10520 16304 10532
rect 15896 10492 16304 10520
rect 15896 10480 15902 10492
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 16850 10520 16856 10532
rect 16540 10492 16856 10520
rect 16540 10480 16546 10492
rect 16850 10480 16856 10492
rect 16908 10480 16914 10532
rect 23109 10523 23167 10529
rect 23109 10489 23121 10523
rect 23155 10520 23167 10523
rect 23155 10492 23428 10520
rect 23155 10489 23167 10492
rect 23109 10483 23167 10489
rect 16206 10452 16212 10464
rect 15028 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 21082 10412 21088 10464
rect 21140 10452 21146 10464
rect 21545 10455 21603 10461
rect 21545 10452 21557 10455
rect 21140 10424 21557 10452
rect 21140 10412 21146 10424
rect 21545 10421 21557 10424
rect 21591 10452 21603 10455
rect 22278 10452 22284 10464
rect 21591 10424 22284 10452
rect 21591 10421 21603 10424
rect 21545 10415 21603 10421
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 23198 10412 23204 10464
rect 23256 10412 23262 10464
rect 23400 10452 23428 10492
rect 24026 10452 24032 10464
rect 23400 10424 24032 10452
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24946 10412 24952 10464
rect 25004 10452 25010 10464
rect 25041 10455 25099 10461
rect 25041 10452 25053 10455
rect 25004 10424 25053 10452
rect 25004 10412 25010 10424
rect 25041 10421 25053 10424
rect 25087 10421 25099 10455
rect 25041 10415 25099 10421
rect 25406 10412 25412 10464
rect 25464 10412 25470 10464
rect 1104 10362 25852 10384
rect 1104 10310 4043 10362
rect 4095 10310 4107 10362
rect 4159 10310 4171 10362
rect 4223 10310 4235 10362
rect 4287 10310 4299 10362
rect 4351 10310 10230 10362
rect 10282 10310 10294 10362
rect 10346 10310 10358 10362
rect 10410 10310 10422 10362
rect 10474 10310 10486 10362
rect 10538 10310 16417 10362
rect 16469 10310 16481 10362
rect 16533 10310 16545 10362
rect 16597 10310 16609 10362
rect 16661 10310 16673 10362
rect 16725 10310 22604 10362
rect 22656 10310 22668 10362
rect 22720 10310 22732 10362
rect 22784 10310 22796 10362
rect 22848 10310 22860 10362
rect 22912 10310 25852 10362
rect 1104 10288 25852 10310
rect 3510 10248 3516 10260
rect 2746 10220 3516 10248
rect 1394 10072 1400 10124
rect 1452 10072 1458 10124
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2746 10112 2774 10220
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 4948 10220 5396 10248
rect 4948 10208 4954 10220
rect 5368 10180 5396 10220
rect 5442 10208 5448 10260
rect 5500 10208 5506 10260
rect 7377 10251 7435 10257
rect 7377 10217 7389 10251
rect 7423 10248 7435 10251
rect 7926 10248 7932 10260
rect 7423 10220 7932 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8478 10248 8484 10260
rect 8435 10220 8484 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 11238 10248 11244 10260
rect 10367 10220 11244 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 12066 10208 12072 10260
rect 12124 10208 12130 10260
rect 13170 10248 13176 10260
rect 12452 10220 13176 10248
rect 6178 10180 6184 10192
rect 5368 10152 6184 10180
rect 6178 10140 6184 10152
rect 6236 10180 6242 10192
rect 10229 10183 10287 10189
rect 6236 10152 7972 10180
rect 6236 10140 6242 10152
rect 1719 10084 2774 10112
rect 5169 10115 5227 10121
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 5169 10081 5181 10115
rect 5215 10112 5227 10115
rect 5902 10112 5908 10124
rect 5215 10084 5908 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 7944 10056 7972 10152
rect 10229 10149 10241 10183
rect 10275 10180 10287 10183
rect 11330 10180 11336 10192
rect 10275 10152 11336 10180
rect 10275 10149 10287 10152
rect 10229 10143 10287 10149
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11974 10140 11980 10192
rect 12032 10140 12038 10192
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10112 9919 10115
rect 11422 10112 11428 10124
rect 9907 10084 11428 10112
rect 9907 10081 9919 10084
rect 9861 10075 9919 10081
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 11606 10072 11612 10124
rect 11664 10072 11670 10124
rect 12452 10121 12480 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 15933 10251 15991 10257
rect 15933 10217 15945 10251
rect 15979 10248 15991 10251
rect 16022 10248 16028 10260
rect 15979 10220 16028 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16669 10251 16727 10257
rect 16669 10217 16681 10251
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 13262 10180 13268 10192
rect 12820 10152 13268 10180
rect 12820 10121 12848 10152
rect 13262 10140 13268 10152
rect 13320 10180 13326 10192
rect 14185 10183 14243 10189
rect 14185 10180 14197 10183
rect 13320 10152 14197 10180
rect 13320 10140 13326 10152
rect 14185 10149 14197 10152
rect 14231 10149 14243 10183
rect 14918 10180 14924 10192
rect 14185 10143 14243 10149
rect 14568 10152 14924 10180
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 13136 10084 13369 10112
rect 13136 10072 13142 10084
rect 13357 10081 13369 10084
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3160 10016 3249 10044
rect 2406 9936 2412 9988
rect 2464 9936 2470 9988
rect 3160 9920 3188 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5092 9976 5120 10007
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5408 10016 5549 10044
rect 5408 10004 5414 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5626 9976 5632 9988
rect 5092 9948 5632 9976
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 3329 9911 3387 9917
rect 3329 9877 3341 9911
rect 3375 9908 3387 9911
rect 3878 9908 3884 9920
rect 3375 9880 3884 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 5736 9908 5764 10007
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 7760 9976 7788 10007
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7984 10016 8033 10044
rect 7984 10004 7990 10016
rect 8021 10013 8033 10016
rect 8067 10044 8079 10047
rect 8202 10044 8208 10056
rect 8067 10016 8208 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8386 10004 8392 10056
rect 8444 10044 8450 10056
rect 8573 10047 8631 10053
rect 8573 10044 8585 10047
rect 8444 10016 8585 10044
rect 8444 10004 8450 10016
rect 8573 10013 8585 10016
rect 8619 10013 8631 10047
rect 8573 10007 8631 10013
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9456 10016 9505 10044
rect 9456 10004 9462 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 10134 10004 10140 10056
rect 10192 10044 10198 10056
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10192 10016 10609 10044
rect 10192 10004 10198 10016
rect 10597 10013 10609 10016
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 11698 10044 11704 10056
rect 11563 10016 11704 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 11348 9976 11376 10007
rect 11698 10004 11704 10016
rect 11756 10044 11762 10056
rect 11882 10044 11888 10056
rect 11756 10016 11888 10044
rect 11756 10004 11762 10016
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12989 10047 13047 10053
rect 12391 10016 12848 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 6972 9948 7972 9976
rect 11348 9948 12434 9976
rect 6972 9936 6978 9948
rect 7944 9920 7972 9948
rect 12406 9920 12434 9948
rect 12618 9936 12624 9988
rect 12676 9936 12682 9988
rect 12710 9936 12716 9988
rect 12768 9936 12774 9988
rect 12820 9976 12848 10016
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13170 10044 13176 10056
rect 13035 10016 13176 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 14568 10053 14596 10152
rect 14918 10140 14924 10152
rect 14976 10180 14982 10192
rect 15013 10183 15071 10189
rect 15013 10180 15025 10183
rect 14976 10152 15025 10180
rect 14976 10140 14982 10152
rect 15013 10149 15025 10152
rect 15059 10149 15071 10183
rect 15562 10180 15568 10192
rect 15013 10143 15071 10149
rect 15120 10152 15568 10180
rect 14734 10072 14740 10124
rect 14792 10072 14798 10124
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 14332 10016 14381 10044
rect 14332 10004 14338 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 15120 10044 15148 10152
rect 15562 10140 15568 10152
rect 15620 10180 15626 10192
rect 16684 10180 16712 10211
rect 16850 10208 16856 10260
rect 16908 10208 16914 10260
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 19886 10248 19892 10260
rect 17184 10220 19892 10248
rect 17184 10208 17190 10220
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20809 10251 20867 10257
rect 20809 10217 20821 10251
rect 20855 10248 20867 10251
rect 22002 10248 22008 10260
rect 20855 10220 22008 10248
rect 20855 10217 20867 10220
rect 20809 10211 20867 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22738 10208 22744 10260
rect 22796 10208 22802 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10248 22891 10251
rect 23014 10248 23020 10260
rect 22879 10220 23020 10248
rect 22879 10217 22891 10220
rect 22833 10211 22891 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23198 10208 23204 10260
rect 23256 10208 23262 10260
rect 25498 10248 25504 10260
rect 23308 10220 25504 10248
rect 15620 10152 16712 10180
rect 15620 10140 15626 10152
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 16482 10112 16488 10124
rect 15243 10084 16488 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 16868 10112 16896 10208
rect 20622 10140 20628 10192
rect 20680 10140 20686 10192
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 22370 10180 22376 10192
rect 21968 10152 22376 10180
rect 21968 10140 21974 10152
rect 22370 10140 22376 10152
rect 22428 10140 22434 10192
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 16868 10084 17325 10112
rect 17313 10081 17325 10084
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10081 19947 10115
rect 19889 10075 19947 10081
rect 14700 10016 15148 10044
rect 14700 10010 14739 10016
rect 14700 10004 14706 10010
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 15654 10004 15660 10056
rect 15712 10004 15718 10056
rect 16040 10053 16436 10054
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10044 15807 10047
rect 16040 10047 16451 10053
rect 16040 10044 16405 10047
rect 15795 10026 16405 10044
rect 15795 10016 16068 10026
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 16393 10013 16405 10026
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 16850 10004 16856 10056
rect 16908 10004 16914 10056
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10013 17095 10047
rect 17037 10007 17095 10013
rect 14645 10001 14703 10004
rect 12894 9976 12900 9988
rect 12820 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9976 12958 9988
rect 13630 9976 13636 9988
rect 12952 9948 13636 9976
rect 12952 9936 12958 9948
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 13725 9979 13783 9985
rect 13725 9945 13737 9979
rect 13771 9976 13783 9979
rect 15194 9976 15200 9988
rect 13771 9948 14596 9976
rect 13771 9945 13783 9948
rect 13725 9939 13783 9945
rect 4856 9880 5764 9908
rect 4856 9868 4862 9880
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 10410 9868 10416 9920
rect 10468 9868 10474 9920
rect 11422 9868 11428 9920
rect 11480 9868 11486 9920
rect 12342 9868 12348 9920
rect 12400 9908 12434 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 12400 9880 13277 9908
rect 12400 9868 12406 9880
rect 13265 9877 13277 9880
rect 13311 9908 13323 9911
rect 14090 9908 14096 9920
rect 13311 9880 14096 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14568 9908 14596 9948
rect 14752 9948 15200 9976
rect 14752 9908 14780 9948
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15304 9976 15332 10004
rect 16025 9979 16083 9985
rect 16025 9976 16037 9979
rect 15304 9948 16037 9976
rect 16025 9945 16037 9948
rect 16071 9945 16083 9979
rect 16025 9939 16083 9945
rect 16207 9979 16265 9985
rect 16207 9945 16219 9979
rect 16253 9945 16265 9979
rect 16207 9939 16265 9945
rect 14568 9880 14780 9908
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 14884 9880 15301 9908
rect 14884 9868 14890 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 15289 9871 15347 9877
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 15838 9908 15844 9920
rect 15712 9880 15844 9908
rect 15712 9868 15718 9880
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16224 9908 16252 9939
rect 16482 9936 16488 9988
rect 16540 9936 16546 9988
rect 16172 9880 16252 9908
rect 16172 9868 16178 9880
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 16868 9917 16896 10004
rect 16685 9911 16743 9917
rect 16685 9908 16697 9911
rect 16448 9880 16697 9908
rect 16448 9868 16454 9880
rect 16685 9877 16697 9880
rect 16731 9877 16743 9911
rect 16685 9871 16743 9877
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9877 16911 9911
rect 17052 9908 17080 10007
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 19610 10004 19616 10056
rect 19668 10004 19674 10056
rect 19904 10044 19932 10075
rect 20346 10072 20352 10124
rect 20404 10072 20410 10124
rect 21358 10112 21364 10124
rect 20456 10084 21364 10112
rect 20456 10044 20484 10084
rect 21358 10072 21364 10084
rect 21416 10112 21422 10124
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 21416 10084 21465 10112
rect 21416 10072 21422 10084
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 19904 10016 20484 10044
rect 20714 10004 20720 10056
rect 20772 10004 20778 10056
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10044 21327 10047
rect 22756 10044 22784 10208
rect 21315 10016 22784 10044
rect 23216 10044 23244 10208
rect 23308 10121 23336 10220
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 23750 10180 23756 10192
rect 23400 10152 23756 10180
rect 23400 10121 23428 10152
rect 23750 10140 23756 10152
rect 23808 10140 23814 10192
rect 24026 10140 24032 10192
rect 24084 10180 24090 10192
rect 24673 10183 24731 10189
rect 24673 10180 24685 10183
rect 24084 10152 24685 10180
rect 24084 10140 24090 10152
rect 24673 10149 24685 10152
rect 24719 10149 24731 10183
rect 24673 10143 24731 10149
rect 23293 10115 23351 10121
rect 23293 10081 23305 10115
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23385 10115 23443 10121
rect 23385 10081 23397 10115
rect 23431 10081 23443 10115
rect 23385 10075 23443 10081
rect 23658 10072 23664 10124
rect 23716 10112 23722 10124
rect 24397 10115 24455 10121
rect 24397 10112 24409 10115
rect 23716 10084 24409 10112
rect 23716 10072 23722 10084
rect 24397 10081 24409 10084
rect 24443 10081 24455 10115
rect 24397 10075 24455 10081
rect 23845 10047 23903 10053
rect 23845 10044 23857 10047
rect 23216 10016 23857 10044
rect 21315 10013 21327 10016
rect 21269 10007 21327 10013
rect 23845 10013 23857 10016
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 24302 10004 24308 10056
rect 24360 10044 24366 10056
rect 25133 10047 25191 10053
rect 25133 10044 25145 10047
rect 24360 10016 25145 10044
rect 24360 10004 24366 10016
rect 25133 10013 25145 10016
rect 25179 10013 25191 10047
rect 25133 10007 25191 10013
rect 20732 9976 20760 10004
rect 21174 9976 21180 9988
rect 20732 9948 21180 9976
rect 21174 9936 21180 9948
rect 21232 9976 21238 9988
rect 21361 9979 21419 9985
rect 21361 9976 21373 9979
rect 21232 9948 21373 9976
rect 21232 9936 21238 9948
rect 21361 9945 21373 9948
rect 21407 9945 21419 9979
rect 21361 9939 21419 9945
rect 21634 9936 21640 9988
rect 21692 9976 21698 9988
rect 23014 9976 23020 9988
rect 21692 9948 23020 9976
rect 21692 9936 21698 9948
rect 23014 9936 23020 9948
rect 23072 9936 23078 9988
rect 17218 9908 17224 9920
rect 17052 9880 17224 9908
rect 16853 9871 16911 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18782 9868 18788 9920
rect 18840 9868 18846 9920
rect 19242 9868 19248 9920
rect 19300 9868 19306 9920
rect 19702 9868 19708 9920
rect 19760 9868 19766 9920
rect 20898 9868 20904 9920
rect 20956 9868 20962 9920
rect 22462 9868 22468 9920
rect 22520 9908 22526 9920
rect 23201 9911 23259 9917
rect 23201 9908 23213 9911
rect 22520 9880 23213 9908
rect 22520 9868 22526 9880
rect 23201 9877 23213 9880
rect 23247 9877 23259 9911
rect 23201 9871 23259 9877
rect 23658 9868 23664 9920
rect 23716 9868 23722 9920
rect 24854 9868 24860 9920
rect 24912 9868 24918 9920
rect 25409 9911 25467 9917
rect 25409 9877 25421 9911
rect 25455 9908 25467 9911
rect 25455 9880 26004 9908
rect 25455 9877 25467 9880
rect 25409 9871 25467 9877
rect 1104 9818 25852 9840
rect 1104 9766 4703 9818
rect 4755 9766 4767 9818
rect 4819 9766 4831 9818
rect 4883 9766 4895 9818
rect 4947 9766 4959 9818
rect 5011 9766 10890 9818
rect 10942 9766 10954 9818
rect 11006 9766 11018 9818
rect 11070 9766 11082 9818
rect 11134 9766 11146 9818
rect 11198 9766 17077 9818
rect 17129 9766 17141 9818
rect 17193 9766 17205 9818
rect 17257 9766 17269 9818
rect 17321 9766 17333 9818
rect 17385 9766 23264 9818
rect 23316 9766 23328 9818
rect 23380 9766 23392 9818
rect 23444 9766 23456 9818
rect 23508 9766 23520 9818
rect 23572 9766 25852 9818
rect 25976 9784 26004 9880
rect 1104 9744 25852 9766
rect 25958 9732 25964 9784
rect 26016 9732 26022 9784
rect 3804 9676 4476 9704
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 3804 9568 3832 9676
rect 4448 9674 4476 9676
rect 4448 9646 4568 9674
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 6270 9704 6276 9716
rect 5500 9676 6276 9704
rect 5500 9664 5506 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 7929 9707 7987 9713
rect 7929 9704 7941 9707
rect 7892 9676 7941 9704
rect 7892 9664 7898 9676
rect 7929 9673 7941 9676
rect 7975 9673 7987 9707
rect 11517 9707 11575 9713
rect 7929 9667 7987 9673
rect 8588 9676 11192 9704
rect 4540 9636 4568 9646
rect 4706 9636 4712 9648
rect 3896 9608 4384 9636
rect 4540 9608 4712 9636
rect 3896 9580 3924 9608
rect 2823 9540 3832 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 1504 9500 1532 9531
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4356 9566 4384 9608
rect 4550 9577 4578 9608
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 5092 9608 5764 9636
rect 5092 9577 5120 9608
rect 5736 9580 5764 9608
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 7616 9608 8064 9636
rect 7616 9596 7622 9608
rect 4433 9571 4491 9577
rect 4433 9566 4445 9571
rect 4356 9538 4445 9566
rect 4433 9537 4445 9538
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5534 9568 5540 9580
rect 5399 9540 5540 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 6086 9528 6092 9580
rect 6144 9528 6150 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7064 9540 7389 9568
rect 7064 9528 7070 9540
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 7742 9568 7748 9580
rect 7423 9540 7748 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 7834 9528 7840 9580
rect 7892 9528 7898 9580
rect 8036 9577 8064 9608
rect 8588 9580 8616 9676
rect 9033 9639 9091 9645
rect 9033 9605 9045 9639
rect 9079 9636 9091 9639
rect 9306 9636 9312 9648
rect 9079 9608 9312 9636
rect 9079 9605 9091 9608
rect 9033 9599 9091 9605
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 10410 9636 10416 9648
rect 10258 9608 10416 9636
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 11164 9580 11192 9676
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11698 9704 11704 9716
rect 11563 9676 11704 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 12158 9704 12164 9716
rect 11848 9676 12164 9704
rect 11848 9664 11854 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 12768 9676 13001 9704
rect 12768 9664 12774 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 13170 9704 13176 9716
rect 12989 9667 13047 9673
rect 13096 9676 13176 9704
rect 12894 9636 12900 9648
rect 11992 9608 12388 9636
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8386 9568 8392 9580
rect 8067 9540 8392 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8570 9528 8576 9580
rect 8628 9528 8634 9580
rect 8754 9528 8760 9580
rect 8812 9528 8818 9580
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11992 9577 12020 9608
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11287 9540 11989 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 12207 9540 12265 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 1504 9472 2697 9500
rect 2685 9469 2697 9472
rect 2731 9500 2743 9503
rect 3142 9500 3148 9512
rect 2731 9472 3148 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 3384 9472 4905 9500
rect 3384 9460 3390 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 5644 9500 5672 9528
rect 6104 9500 6132 9528
rect 11054 9500 11060 9512
rect 5215 9472 5672 9500
rect 5736 9472 6132 9500
rect 7944 9472 11060 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 5261 9435 5319 9441
rect 3651 9404 4660 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 992 9336 1593 9364
rect 992 9324 998 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3142 9364 3148 9376
rect 3099 9336 3148 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3142 9324 3148 9336
rect 3200 9364 3206 9376
rect 3620 9364 3648 9395
rect 4632 9376 4660 9404
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5736 9432 5764 9472
rect 5307 9404 5764 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 7944 9376 7972 9472
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11882 9460 11888 9512
rect 11940 9460 11946 9512
rect 12360 9500 12388 9608
rect 12452 9608 12900 9636
rect 12452 9577 12480 9608
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 13096 9645 13124 9676
rect 13170 9664 13176 9676
rect 13228 9704 13234 9716
rect 13228 9676 13860 9704
rect 13228 9664 13234 9676
rect 13081 9639 13139 9645
rect 13081 9605 13093 9639
rect 13127 9636 13139 9639
rect 13127 9608 13161 9636
rect 13127 9605 13139 9608
rect 13081 9599 13139 9605
rect 13262 9596 13268 9648
rect 13320 9645 13326 9648
rect 13320 9639 13339 9645
rect 13327 9605 13339 9639
rect 13725 9639 13783 9645
rect 13725 9636 13737 9639
rect 13320 9599 13339 9605
rect 13372 9608 13737 9636
rect 13320 9596 13326 9599
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12526 9528 12532 9580
rect 12584 9577 12590 9580
rect 12584 9568 12596 9577
rect 12805 9571 12863 9577
rect 12805 9570 12817 9571
rect 12584 9540 12629 9568
rect 12728 9542 12817 9570
rect 12584 9531 12596 9540
rect 12584 9528 12590 9531
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 12360 9472 12633 9500
rect 12621 9469 12633 9472
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 10134 9392 10140 9444
rect 10192 9392 10198 9444
rect 11900 9432 11928 9460
rect 12728 9432 12756 9542
rect 12805 9537 12817 9542
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 11900 9404 12756 9432
rect 3200 9336 3648 9364
rect 3200 9324 3206 9336
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3752 9336 3801 9364
rect 3752 9324 3758 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9364 4031 9367
rect 4430 9364 4436 9376
rect 4019 9336 4436 9364
rect 4019 9333 4031 9336
rect 3973 9327 4031 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 7653 9367 7711 9373
rect 7653 9333 7665 9367
rect 7699 9364 7711 9367
rect 7926 9364 7932 9376
rect 7699 9336 7932 9364
rect 7699 9333 7711 9336
rect 7653 9327 7711 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10152 9364 10180 9392
rect 9824 9336 10180 9364
rect 10505 9367 10563 9373
rect 9824 9324 9830 9336
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 10686 9364 10692 9376
rect 10551 9336 10692 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13136 9336 13277 9364
rect 13136 9324 13142 9336
rect 13265 9333 13277 9336
rect 13311 9364 13323 9367
rect 13372 9364 13400 9608
rect 13725 9605 13737 9608
rect 13771 9605 13783 9639
rect 13832 9636 13860 9676
rect 17494 9664 17500 9716
rect 17552 9664 17558 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18104 9676 18276 9704
rect 18104 9664 18110 9676
rect 14737 9639 14795 9645
rect 14737 9636 14749 9639
rect 13832 9608 14749 9636
rect 13725 9599 13783 9605
rect 14737 9605 14749 9608
rect 14783 9605 14795 9639
rect 14737 9599 14795 9605
rect 15028 9608 15332 9636
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13688 9540 13921 9568
rect 13688 9528 13694 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14016 9500 14044 9531
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 15028 9577 15056 9608
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 15013 9571 15071 9577
rect 14691 9540 14872 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14844 9512 14872 9540
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15304 9568 15332 9608
rect 15378 9596 15384 9648
rect 15436 9596 15442 9648
rect 15580 9608 16528 9636
rect 15580 9577 15608 9608
rect 16500 9580 16528 9608
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15304 9540 15577 9568
rect 15197 9531 15255 9537
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 13464 9472 14044 9500
rect 13464 9441 13492 9472
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14332 9472 14780 9500
rect 14332 9460 14338 9472
rect 13449 9435 13507 9441
rect 13449 9401 13461 9435
rect 13495 9401 13507 9435
rect 14752 9432 14780 9472
rect 14826 9460 14832 9512
rect 14884 9460 14890 9512
rect 15212 9500 15240 9531
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 15712 9540 15761 9568
rect 15712 9528 15718 9540
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9537 15991 9571
rect 15933 9531 15991 9537
rect 15286 9500 15292 9512
rect 15212 9472 15292 9500
rect 15286 9460 15292 9472
rect 15344 9500 15350 9512
rect 15948 9500 15976 9531
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 16080 9540 16129 9568
rect 16080 9528 16086 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 17512 9568 17540 9664
rect 18248 9580 18276 9676
rect 19996 9676 22094 9704
rect 19794 9596 19800 9648
rect 19852 9636 19858 9648
rect 19996 9645 20024 9676
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 19852 9608 19993 9636
rect 19852 9596 19858 9608
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 22066 9636 22094 9676
rect 23106 9664 23112 9716
rect 23164 9664 23170 9716
rect 23750 9664 23756 9716
rect 23808 9704 23814 9716
rect 23808 9676 24256 9704
rect 23808 9664 23814 9676
rect 23124 9636 23152 9664
rect 22066 9608 23152 9636
rect 19981 9599 20039 9605
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 17512 9540 17601 9568
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 22664 9577 22692 9608
rect 23658 9596 23664 9648
rect 23716 9596 23722 9648
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 20864 9540 21465 9568
rect 20864 9528 20870 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 15344 9472 15976 9500
rect 15344 9460 15350 9472
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16632 9472 16773 9500
rect 16632 9460 16638 9472
rect 16761 9469 16773 9472
rect 16807 9500 16819 9503
rect 18782 9500 18788 9512
rect 16807 9472 18788 9500
rect 16807 9469 16819 9472
rect 16761 9463 16819 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 22922 9460 22928 9512
rect 22980 9460 22986 9512
rect 24228 9500 24256 9676
rect 24854 9664 24860 9716
rect 24912 9664 24918 9716
rect 24946 9664 24952 9716
rect 25004 9664 25010 9716
rect 24872 9636 24900 9664
rect 24872 9608 25544 9636
rect 24854 9528 24860 9580
rect 24912 9528 24918 9580
rect 25516 9577 25544 9608
rect 25501 9571 25559 9577
rect 25501 9537 25513 9571
rect 25547 9537 25559 9571
rect 25501 9531 25559 9537
rect 24762 9500 24768 9512
rect 24228 9472 24768 9500
rect 24762 9460 24768 9472
rect 24820 9500 24826 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 24820 9472 25053 9500
rect 24820 9460 24826 9472
rect 25041 9469 25053 9472
rect 25087 9469 25099 9503
rect 25041 9463 25099 9469
rect 15470 9432 15476 9444
rect 14752 9404 15476 9432
rect 13449 9395 13507 9401
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 16025 9435 16083 9441
rect 16025 9432 16037 9435
rect 15896 9404 16037 9432
rect 15896 9392 15902 9404
rect 16025 9401 16037 9404
rect 16071 9432 16083 9435
rect 16666 9432 16672 9444
rect 16071 9404 16672 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17034 9392 17040 9444
rect 17092 9432 17098 9444
rect 24397 9435 24455 9441
rect 17092 9404 22094 9432
rect 17092 9392 17098 9404
rect 13311 9336 13400 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 15160 9336 17325 9364
rect 15160 9324 15166 9336
rect 17313 9333 17325 9336
rect 17359 9333 17371 9367
rect 17313 9327 17371 9333
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 18322 9364 18328 9376
rect 17911 9336 18328 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 21266 9324 21272 9376
rect 21324 9324 21330 9376
rect 22066 9364 22094 9404
rect 24397 9401 24409 9435
rect 24443 9401 24455 9435
rect 24397 9395 24455 9401
rect 24412 9364 24440 9395
rect 22066 9336 24440 9364
rect 24486 9324 24492 9376
rect 24544 9324 24550 9376
rect 25314 9324 25320 9376
rect 25372 9324 25378 9376
rect 1104 9274 25852 9296
rect 1104 9222 4043 9274
rect 4095 9222 4107 9274
rect 4159 9222 4171 9274
rect 4223 9222 4235 9274
rect 4287 9222 4299 9274
rect 4351 9222 10230 9274
rect 10282 9222 10294 9274
rect 10346 9222 10358 9274
rect 10410 9222 10422 9274
rect 10474 9222 10486 9274
rect 10538 9222 16417 9274
rect 16469 9222 16481 9274
rect 16533 9222 16545 9274
rect 16597 9222 16609 9274
rect 16661 9222 16673 9274
rect 16725 9222 22604 9274
rect 22656 9222 22668 9274
rect 22720 9222 22732 9274
rect 22784 9222 22796 9274
rect 22848 9222 22860 9274
rect 22912 9222 25852 9274
rect 1104 9200 25852 9222
rect 3142 9120 3148 9172
rect 3200 9120 3206 9172
rect 3326 9120 3332 9172
rect 3384 9120 3390 9172
rect 3436 9132 5672 9160
rect 3160 8965 3188 9120
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 3344 9024 3372 9120
rect 3283 8996 3372 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3436 8968 3464 9132
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4706 9092 4712 9104
rect 4212 9064 4712 9092
rect 4212 9052 4218 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 5534 9092 5540 9104
rect 4908 9064 5540 9092
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 3559 8996 4261 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4338 8984 4344 9036
rect 4396 8984 4402 9036
rect 4430 8984 4436 9036
rect 4488 8984 4494 9036
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 4580 8996 4844 9024
rect 4580 8984 4586 8996
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3936 8928 4169 8956
rect 3936 8916 3942 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4448 8956 4476 8984
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4448 8928 4721 8956
rect 4157 8919 4215 8925
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4816 8888 4844 8996
rect 4908 8965 4936 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 5644 9092 5672 9132
rect 5718 9120 5724 9172
rect 5776 9120 5782 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9677 9163 9735 9169
rect 8352 9132 9536 9160
rect 8352 9120 8358 9132
rect 8570 9092 8576 9104
rect 5644 9064 8576 9092
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 9508 9101 9536 9132
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9766 9160 9772 9172
rect 9723 9132 9772 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10060 9132 12664 9160
rect 9493 9095 9551 9101
rect 9493 9061 9505 9095
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 10060 9092 10088 9132
rect 9640 9064 10088 9092
rect 9640 9052 9646 9064
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5350 9024 5356 9036
rect 5031 8996 5356 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5350 8984 5356 8996
rect 5408 9024 5414 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5408 8996 5641 9024
rect 5408 8984 5414 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 8662 9024 8668 9036
rect 6328 8996 8668 9024
rect 6328 8984 6334 8996
rect 8662 8984 8668 8996
rect 8720 9024 8726 9036
rect 9784 9033 9812 9064
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 11756 9064 12265 9092
rect 11756 9052 11762 9064
rect 12253 9061 12265 9064
rect 12299 9061 12311 9095
rect 12253 9055 12311 9061
rect 12342 9052 12348 9104
rect 12400 9052 12406 9104
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8720 8996 9229 9024
rect 8720 8984 8726 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 11204 8996 11437 9024
rect 11204 8984 11210 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5092 8888 5120 8919
rect 4816 8860 5120 8888
rect 5276 8888 5304 8919
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9364 8950 9720 8956
rect 9784 8950 9965 8956
rect 9364 8928 9965 8950
rect 9364 8916 9370 8928
rect 9692 8922 9812 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 5828 8888 5856 8916
rect 5276 8860 5856 8888
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 5276 8820 5304 8860
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 11238 8888 11244 8900
rect 8260 8860 11244 8888
rect 8260 8848 8266 8860
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 11440 8888 11468 8987
rect 11882 8984 11888 9036
rect 11940 8984 11946 9036
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12636 9024 12664 9132
rect 13170 9120 13176 9172
rect 13228 9120 13234 9172
rect 14182 9120 14188 9172
rect 14240 9120 14246 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 16022 9160 16028 9172
rect 14884 9132 16028 9160
rect 14884 9120 14890 9132
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19686 9163 19744 9169
rect 19686 9160 19698 9163
rect 18923 9132 19698 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19686 9129 19698 9132
rect 19732 9129 19744 9163
rect 19686 9123 19744 9129
rect 20898 9120 20904 9172
rect 20956 9120 20962 9172
rect 21174 9120 21180 9172
rect 21232 9120 21238 9172
rect 22922 9120 22928 9172
rect 22980 9160 22986 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 22980 9132 23305 9160
rect 22980 9120 22986 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 24486 9120 24492 9172
rect 24544 9160 24550 9172
rect 24544 9132 25360 9160
rect 24544 9120 24550 9132
rect 13188 9092 13216 9120
rect 13998 9092 14004 9104
rect 13188 9064 14004 9092
rect 12894 9024 12900 9036
rect 12636 8996 12900 9024
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 11992 8956 12020 8984
rect 12636 8965 12664 8996
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13188 9024 13216 9064
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 14200 9024 14228 9120
rect 15194 9052 15200 9104
rect 15252 9052 15258 9104
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 17678 9092 17684 9104
rect 16908 9064 17684 9092
rect 16908 9052 16914 9064
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 13096 8996 13216 9024
rect 13280 8996 14228 9024
rect 15212 9024 15240 9052
rect 18690 9024 18696 9036
rect 15212 8996 18696 9024
rect 13096 8965 13124 8996
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11563 8928 12173 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8925 12679 8959
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12621 8919 12679 8925
rect 12912 8928 13001 8956
rect 12452 8888 12480 8919
rect 12912 8888 12940 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13280 8956 13308 8996
rect 18690 8984 18696 8996
rect 18748 8984 18754 9036
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19794 9024 19800 9036
rect 19475 8996 19800 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 20916 9024 20944 9120
rect 23676 9064 25268 9092
rect 23676 9033 23704 9064
rect 25240 9036 25268 9064
rect 23661 9027 23719 9033
rect 20916 8996 21496 9024
rect 13219 8928 13308 8956
rect 13357 8959 13415 8965
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13538 8956 13544 8968
rect 13403 8928 13544 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13538 8916 13544 8928
rect 13596 8956 13602 8968
rect 14458 8956 14464 8968
rect 13596 8928 14464 8956
rect 13596 8916 13602 8928
rect 14458 8916 14464 8928
rect 14516 8956 14522 8968
rect 16022 8956 16028 8968
rect 14516 8928 16028 8956
rect 14516 8916 14522 8928
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16206 8916 16212 8968
rect 16264 8916 16270 8968
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 17034 8956 17040 8968
rect 16724 8928 17040 8956
rect 16724 8916 16730 8928
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18012 8928 18245 8956
rect 18012 8916 18018 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8956 19119 8959
rect 19242 8956 19248 8968
rect 19107 8928 19248 8956
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 21266 8956 21272 8968
rect 20838 8928 21272 8956
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 21468 8965 21496 8996
rect 23661 8993 23673 9027
rect 23707 8993 23719 9027
rect 23661 8987 23719 8993
rect 24762 8984 24768 9036
rect 24820 9024 24826 9036
rect 24949 9027 25007 9033
rect 24949 9024 24961 9027
rect 24820 8996 24961 9024
rect 24820 8984 24826 8996
rect 24949 8993 24961 8996
rect 24995 8993 25007 9027
rect 24949 8987 25007 8993
rect 25222 8984 25228 9036
rect 25280 8984 25286 9036
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8925 23535 8959
rect 25332 8956 25360 9132
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25332 8928 25513 8956
rect 23477 8919 23535 8925
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 15102 8888 15108 8900
rect 11440 8860 12848 8888
rect 12912 8860 15108 8888
rect 4488 8792 5304 8820
rect 5445 8823 5503 8829
rect 4488 8780 4494 8792
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 5810 8820 5816 8832
rect 5491 8792 5816 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 5902 8780 5908 8832
rect 5960 8780 5966 8832
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 9456 8792 10149 8820
rect 9456 8780 9462 8792
rect 10137 8789 10149 8792
rect 10183 8789 10195 8823
rect 10137 8783 10195 8789
rect 11974 8780 11980 8832
rect 12032 8780 12038 8832
rect 12710 8780 12716 8832
rect 12768 8780 12774 8832
rect 12820 8820 12848 8860
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 15654 8848 15660 8900
rect 15712 8888 15718 8900
rect 15712 8860 18184 8888
rect 15712 8848 15718 8860
rect 14182 8820 14188 8832
rect 12820 8792 14188 8820
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 16758 8780 16764 8832
rect 16816 8780 16822 8832
rect 17494 8780 17500 8832
rect 17552 8780 17558 8832
rect 18046 8780 18052 8832
rect 18104 8780 18110 8832
rect 18156 8820 18184 8860
rect 21008 8860 22048 8888
rect 21008 8820 21036 8860
rect 22020 8832 22048 8860
rect 18156 8792 21036 8820
rect 21266 8780 21272 8832
rect 21324 8780 21330 8832
rect 22002 8780 22008 8832
rect 22060 8780 22066 8832
rect 23492 8820 23520 8919
rect 24213 8891 24271 8897
rect 24213 8857 24225 8891
rect 24259 8888 24271 8891
rect 24857 8891 24915 8897
rect 24857 8888 24869 8891
rect 24259 8860 24869 8888
rect 24259 8857 24271 8860
rect 24213 8851 24271 8857
rect 24857 8857 24869 8860
rect 24903 8857 24915 8891
rect 24857 8851 24915 8857
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 23492 8792 24409 8820
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 24397 8783 24455 8789
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 25317 8823 25375 8829
rect 25317 8789 25329 8823
rect 25363 8820 25375 8823
rect 25363 8792 25912 8820
rect 25363 8789 25375 8792
rect 25317 8783 25375 8789
rect 1104 8730 25852 8752
rect 1104 8678 4703 8730
rect 4755 8678 4767 8730
rect 4819 8678 4831 8730
rect 4883 8678 4895 8730
rect 4947 8678 4959 8730
rect 5011 8678 10890 8730
rect 10942 8678 10954 8730
rect 11006 8678 11018 8730
rect 11070 8678 11082 8730
rect 11134 8678 11146 8730
rect 11198 8678 17077 8730
rect 17129 8678 17141 8730
rect 17193 8678 17205 8730
rect 17257 8678 17269 8730
rect 17321 8678 17333 8730
rect 17385 8678 23264 8730
rect 23316 8678 23328 8730
rect 23380 8678 23392 8730
rect 23444 8678 23456 8730
rect 23508 8678 23520 8730
rect 23572 8678 25852 8730
rect 1104 8656 25852 8678
rect 3786 8616 3792 8628
rect 2746 8588 3792 8616
rect 2746 8548 2774 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 5350 8576 5356 8628
rect 5408 8576 5414 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 9306 8576 9312 8628
rect 9364 8576 9370 8628
rect 12618 8616 12624 8628
rect 11256 8588 12624 8616
rect 1964 8520 2774 8548
rect 1964 8489 1992 8520
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8449 1547 8483
rect 1489 8443 1547 8449
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 1504 8412 1532 8443
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 2096 8452 2145 8480
rect 2096 8440 2102 8452
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 3694 8440 3700 8492
rect 3752 8489 3758 8492
rect 3752 8480 3764 8489
rect 3752 8452 3797 8480
rect 3752 8443 3764 8452
rect 3752 8440 3758 8443
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3936 8452 3985 8480
rect 3936 8440 3942 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4672 8452 4905 8480
rect 4672 8440 4678 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 3418 8412 3424 8424
rect 1504 8384 3424 8412
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 4706 8412 4712 8424
rect 4571 8384 4712 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 7852 8412 7880 8576
rect 9674 8508 9680 8560
rect 9732 8508 9738 8560
rect 9766 8508 9772 8560
rect 9824 8508 9830 8560
rect 10778 8548 10784 8560
rect 9876 8520 10784 8548
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 9582 8480 9588 8492
rect 8444 8452 9588 8480
rect 8444 8440 8450 8452
rect 9582 8440 9588 8452
rect 9640 8480 9646 8492
rect 9876 8480 9904 8520
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 9640 8452 9904 8480
rect 9640 8440 9646 8452
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 7791 8384 7880 8412
rect 9646 8384 9965 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 1670 8304 1676 8356
rect 1728 8304 1734 8356
rect 2317 8347 2375 8353
rect 2317 8313 2329 8347
rect 2363 8344 2375 8347
rect 2774 8344 2780 8356
rect 2363 8316 2780 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 9646 8344 9674 8384
rect 9953 8381 9965 8384
rect 9999 8412 10011 8415
rect 11256 8412 11284 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 12952 8588 14044 8616
rect 12952 8576 12958 8588
rect 11440 8520 12112 8548
rect 11440 8492 11468 8520
rect 11422 8440 11428 8492
rect 11480 8440 11486 8492
rect 11885 8484 11943 8489
rect 11974 8484 11980 8492
rect 11885 8483 11980 8484
rect 11885 8449 11897 8483
rect 11931 8456 11980 8483
rect 11931 8449 11943 8456
rect 11885 8443 11943 8449
rect 11974 8440 11980 8456
rect 12032 8440 12038 8492
rect 12084 8489 12112 8520
rect 12250 8508 12256 8560
rect 12308 8508 12314 8560
rect 12710 8508 12716 8560
rect 12768 8508 12774 8560
rect 14016 8548 14044 8588
rect 14182 8576 14188 8628
rect 14240 8576 14246 8628
rect 15654 8576 15660 8628
rect 15712 8576 15718 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16758 8616 16764 8628
rect 15795 8588 16764 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17129 8619 17187 8625
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17678 8616 17684 8628
rect 17175 8588 17684 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18138 8616 18144 8628
rect 17880 8588 18144 8616
rect 17880 8548 17908 8588
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19944 8588 19993 8616
rect 19944 8576 19950 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 19981 8579 20039 8585
rect 20806 8576 20812 8628
rect 20864 8576 20870 8628
rect 21453 8619 21511 8625
rect 21453 8585 21465 8619
rect 21499 8585 21511 8619
rect 25884 8616 25912 8792
rect 21453 8579 21511 8585
rect 24044 8588 25912 8616
rect 14016 8520 15976 8548
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 12268 8480 12296 8508
rect 12207 8452 12296 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15243 8452 15332 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 9999 8384 11284 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 12250 8372 12256 8424
rect 12308 8412 12314 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12308 8384 12449 8412
rect 12308 8372 12314 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 4396 8316 9674 8344
rect 4396 8304 4402 8316
rect 11698 8304 11704 8356
rect 11756 8304 11762 8356
rect 15304 8353 15332 8452
rect 15948 8421 15976 8520
rect 16960 8520 17908 8548
rect 16960 8489 16988 8520
rect 18046 8508 18052 8560
rect 18104 8508 18110 8560
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 20993 8551 21051 8557
rect 20993 8548 21005 8551
rect 20404 8520 21005 8548
rect 20404 8508 20410 8520
rect 20993 8517 21005 8520
rect 21039 8517 21051 8551
rect 20993 8511 21051 8517
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8449 19947 8483
rect 21468 8480 21496 8579
rect 24044 8557 24072 8588
rect 24029 8551 24087 8557
rect 24029 8517 24041 8551
rect 24075 8517 24087 8551
rect 25314 8548 25320 8560
rect 25254 8520 25320 8548
rect 24029 8511 24087 8517
rect 25314 8508 25320 8520
rect 25372 8508 25378 8560
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21468 8452 22017 8480
rect 19889 8443 19947 8449
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 15979 8384 16773 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 17218 8372 17224 8424
rect 17276 8372 17282 8424
rect 17494 8372 17500 8424
rect 17552 8372 17558 8424
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 19904 8412 19932 8443
rect 18748 8384 19932 8412
rect 18748 8372 18754 8384
rect 20714 8372 20720 8424
rect 20772 8372 20778 8424
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 21100 8384 23765 8412
rect 15289 8347 15347 8353
rect 15289 8313 15301 8347
rect 15335 8313 15347 8347
rect 15289 8307 15347 8313
rect 20622 8304 20628 8356
rect 20680 8304 20686 8356
rect 20732 8344 20760 8372
rect 21100 8344 21128 8384
rect 23753 8381 23765 8384
rect 23799 8381 23811 8415
rect 23753 8375 23811 8381
rect 23860 8384 25912 8412
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 20732 8316 21128 8344
rect 21192 8316 21281 8344
rect 1946 8236 1952 8288
rect 2004 8236 2010 8288
rect 3510 8236 3516 8288
rect 3568 8236 3574 8288
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4856 8248 4997 8276
rect 4856 8236 4862 8248
rect 4985 8245 4997 8248
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 12158 8276 12164 8288
rect 7892 8248 12164 8276
rect 7892 8236 7898 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 15010 8236 15016 8288
rect 15068 8236 15074 8288
rect 18046 8236 18052 8288
rect 18104 8276 18110 8288
rect 18969 8279 19027 8285
rect 18969 8276 18981 8279
rect 18104 8248 18981 8276
rect 18104 8236 18110 8248
rect 18969 8245 18981 8248
rect 19015 8245 19027 8279
rect 20640 8276 20668 8304
rect 21192 8276 21220 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21821 8347 21879 8353
rect 21821 8313 21833 8347
rect 21867 8344 21879 8347
rect 21867 8316 21956 8344
rect 21867 8313 21879 8316
rect 21821 8307 21879 8313
rect 20640 8248 21220 8276
rect 21928 8276 21956 8316
rect 22002 8304 22008 8356
rect 22060 8344 22066 8356
rect 23860 8344 23888 8384
rect 25884 8356 25912 8384
rect 22060 8316 23888 8344
rect 22060 8304 22066 8316
rect 25222 8304 25228 8356
rect 25280 8344 25286 8356
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 25280 8316 25513 8344
rect 25280 8304 25286 8316
rect 25501 8313 25513 8316
rect 25547 8313 25559 8347
rect 25501 8307 25559 8313
rect 25866 8304 25872 8356
rect 25924 8304 25930 8356
rect 22094 8276 22100 8288
rect 21928 8248 22100 8276
rect 18969 8239 19027 8245
rect 22094 8236 22100 8248
rect 22152 8236 22158 8288
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 23106 8276 23112 8288
rect 22244 8248 23112 8276
rect 22244 8236 22250 8248
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 1104 8186 25852 8208
rect 1104 8134 4043 8186
rect 4095 8134 4107 8186
rect 4159 8134 4171 8186
rect 4223 8134 4235 8186
rect 4287 8134 4299 8186
rect 4351 8134 10230 8186
rect 10282 8134 10294 8186
rect 10346 8134 10358 8186
rect 10410 8134 10422 8186
rect 10474 8134 10486 8186
rect 10538 8134 16417 8186
rect 16469 8134 16481 8186
rect 16533 8134 16545 8186
rect 16597 8134 16609 8186
rect 16661 8134 16673 8186
rect 16725 8134 22604 8186
rect 22656 8134 22668 8186
rect 22720 8134 22732 8186
rect 22784 8134 22796 8186
rect 22848 8134 22860 8186
rect 22912 8134 25852 8186
rect 1104 8112 25852 8134
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 3844 8044 4261 8072
rect 3844 8032 3850 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 7374 8032 7380 8084
rect 7432 8032 7438 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7708 8044 7941 8072
rect 7708 8032 7714 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8754 8072 8760 8084
rect 8343 8044 8760 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9766 8072 9772 8084
rect 9539 8044 9772 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 13814 8072 13820 8084
rect 13771 8044 13820 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 13906 8032 13912 8084
rect 13964 8032 13970 8084
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 16264 8044 16405 8072
rect 16264 8032 16270 8044
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 17954 8032 17960 8084
rect 18012 8032 18018 8084
rect 18138 8032 18144 8084
rect 18196 8032 18202 8084
rect 18414 8032 18420 8084
rect 18472 8032 18478 8084
rect 4430 8004 4436 8016
rect 2746 7976 4436 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 2746 7936 2774 7976
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 6086 7964 6092 8016
rect 6144 8004 6150 8016
rect 7392 8004 7420 8032
rect 8202 8004 8208 8016
rect 6144 7976 7328 8004
rect 7392 7976 8208 8004
rect 6144 7964 6150 7976
rect 1443 7908 2774 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 3881 7939 3939 7945
rect 3881 7936 3893 7939
rect 3568 7908 3893 7936
rect 3568 7896 3574 7908
rect 3881 7905 3893 7908
rect 3927 7905 3939 7939
rect 4798 7936 4804 7948
rect 3881 7899 3939 7905
rect 3988 7908 4804 7936
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 3988 7877 4016 7908
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6914 7936 6920 7948
rect 5868 7908 6920 7936
rect 5868 7896 5874 7908
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 6972 7908 7052 7936
rect 6972 7896 6978 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4614 7868 4620 7880
rect 4571 7840 4620 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 1946 7800 1952 7812
rect 1719 7772 1952 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 1946 7760 1952 7772
rect 2004 7760 2010 7812
rect 4448 7800 4476 7831
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6546 7868 6552 7880
rect 5960 7840 6552 7868
rect 5960 7828 5966 7840
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 7024 7877 7052 7908
rect 7009 7871 7067 7877
rect 6656 7840 6960 7868
rect 4706 7800 4712 7812
rect 3160 7772 4712 7800
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3160 7741 3188 7772
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 6086 7760 6092 7812
rect 6144 7800 6150 7812
rect 6365 7803 6423 7809
rect 6365 7800 6377 7803
rect 6144 7772 6377 7800
rect 6144 7760 6150 7772
rect 6365 7769 6377 7772
rect 6411 7769 6423 7803
rect 6365 7763 6423 7769
rect 3145 7735 3203 7741
rect 3145 7732 3157 7735
rect 3108 7704 3157 7732
rect 3108 7692 3114 7704
rect 3145 7701 3157 7704
rect 3191 7701 3203 7735
rect 3145 7695 3203 7701
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 6656 7732 6684 7840
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 6932 7800 6960 7840
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7300 7868 7328 7976
rect 8202 7964 8208 7976
rect 8260 8004 8266 8016
rect 8481 8007 8539 8013
rect 8481 8004 8493 8007
rect 8260 7976 8493 8004
rect 8260 7964 8266 7976
rect 8481 7973 8493 7976
rect 8527 7973 8539 8007
rect 8481 7967 8539 7973
rect 8662 7964 8668 8016
rect 8720 7964 8726 8016
rect 11238 7964 11244 8016
rect 11296 8004 11302 8016
rect 12250 8004 12256 8016
rect 11296 7976 12256 8004
rect 11296 7964 11302 7976
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 13354 7964 13360 8016
rect 13412 8004 13418 8016
rect 13449 8007 13507 8013
rect 13449 8004 13461 8007
rect 13412 7976 13461 8004
rect 13412 7964 13418 7976
rect 13449 7973 13461 7976
rect 13495 7973 13507 8007
rect 13924 8004 13952 8032
rect 13449 7967 13507 7973
rect 13556 7976 14596 8004
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 7466 7936 7472 7948
rect 7423 7908 7472 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8352 7908 9045 7936
rect 8352 7896 8358 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13556 7936 13584 7976
rect 13219 7908 13584 7936
rect 13633 7939 13691 7945
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 13679 7908 13952 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 7742 7868 7748 7880
rect 7300 7840 7748 7868
rect 7009 7831 7067 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8478 7868 8484 7880
rect 8067 7840 8484 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8846 7868 8852 7880
rect 8619 7840 8852 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 13924 7877 13952 7908
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 11882 7800 11888 7812
rect 6932 7772 11888 7800
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 3660 7704 6684 7732
rect 6733 7735 6791 7741
rect 3660 7692 3666 7704
rect 6733 7701 6745 7735
rect 6779 7732 6791 7735
rect 7098 7732 7104 7744
rect 6779 7704 7104 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8938 7732 8944 7744
rect 8260 7704 8944 7732
rect 8260 7692 8266 7704
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 14182 7732 14188 7744
rect 11664 7704 14188 7732
rect 11664 7692 11670 7704
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14568 7732 14596 7976
rect 17494 7964 17500 8016
rect 17552 8004 17558 8016
rect 17770 8004 17776 8016
rect 17552 7976 17776 8004
rect 17552 7964 17558 7976
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7936 14703 7939
rect 17218 7936 17224 7948
rect 14691 7908 17224 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 17218 7896 17224 7908
rect 17276 7936 17282 7948
rect 17276 7908 17908 7936
rect 17276 7896 17282 7908
rect 17880 7880 17908 7908
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16632 7840 17816 7868
rect 16632 7828 16638 7840
rect 17788 7812 17816 7840
rect 17862 7828 17868 7880
rect 17920 7828 17926 7880
rect 18432 7868 18460 8032
rect 22186 7964 22192 8016
rect 22244 8004 22250 8016
rect 25317 8007 25375 8013
rect 25317 8004 25329 8007
rect 22244 7976 25329 8004
rect 22244 7964 22250 7976
rect 25317 7973 25329 7976
rect 25363 7973 25375 8007
rect 25317 7967 25375 7973
rect 18690 7896 18696 7948
rect 18748 7896 18754 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21174 7936 21180 7948
rect 21131 7908 21180 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 17972 7840 18460 7868
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7800 14979 7803
rect 15010 7800 15016 7812
rect 14967 7772 15016 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 15562 7760 15568 7812
rect 15620 7760 15626 7812
rect 17497 7803 17555 7809
rect 17497 7769 17509 7803
rect 17543 7769 17555 7803
rect 17497 7763 17555 7769
rect 17512 7732 17540 7763
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 17972 7800 18000 7840
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 20772 7840 20821 7868
rect 20772 7828 20778 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 25041 7871 25099 7877
rect 22152 7840 22218 7868
rect 22152 7828 22158 7840
rect 25041 7837 25053 7871
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 25958 7868 25964 7880
rect 25547 7840 25964 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 17828 7772 18000 7800
rect 17828 7760 17834 7772
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 18601 7803 18659 7809
rect 18601 7800 18613 7803
rect 18472 7772 18613 7800
rect 18472 7760 18478 7772
rect 18601 7769 18613 7772
rect 18647 7769 18659 7803
rect 25056 7800 25084 7831
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 25056 7772 25728 7800
rect 18601 7763 18659 7769
rect 25700 7744 25728 7772
rect 17678 7732 17684 7744
rect 14568 7704 17684 7732
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 19242 7732 19248 7744
rect 18555 7704 19248 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22557 7735 22615 7741
rect 22557 7732 22569 7735
rect 22152 7704 22569 7732
rect 22152 7692 22158 7704
rect 22557 7701 22569 7704
rect 22603 7701 22615 7735
rect 22557 7695 22615 7701
rect 24946 7692 24952 7744
rect 25004 7732 25010 7744
rect 25225 7735 25283 7741
rect 25225 7732 25237 7735
rect 25004 7704 25237 7732
rect 25004 7692 25010 7704
rect 25225 7701 25237 7704
rect 25271 7701 25283 7735
rect 25225 7695 25283 7701
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 1104 7642 25852 7664
rect 1104 7590 4703 7642
rect 4755 7590 4767 7642
rect 4819 7590 4831 7642
rect 4883 7590 4895 7642
rect 4947 7590 4959 7642
rect 5011 7590 10890 7642
rect 10942 7590 10954 7642
rect 11006 7590 11018 7642
rect 11070 7590 11082 7642
rect 11134 7590 11146 7642
rect 11198 7590 17077 7642
rect 17129 7590 17141 7642
rect 17193 7590 17205 7642
rect 17257 7590 17269 7642
rect 17321 7590 17333 7642
rect 17385 7590 23264 7642
rect 23316 7590 23328 7642
rect 23380 7590 23392 7642
rect 23444 7590 23456 7642
rect 23508 7590 23520 7642
rect 23572 7590 25852 7642
rect 1104 7568 25852 7590
rect 934 7488 940 7540
rect 992 7528 998 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 992 7500 1593 7528
rect 992 7488 998 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 7098 7528 7104 7540
rect 5920 7500 7104 7528
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7460 1547 7463
rect 2038 7460 2044 7472
rect 1535 7432 2044 7460
rect 1535 7429 1547 7432
rect 1489 7423 1547 7429
rect 2038 7420 2044 7432
rect 2096 7420 2102 7472
rect 5920 7469 5948 7500
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7282 7488 7288 7540
rect 7340 7488 7346 7540
rect 8386 7528 8392 7540
rect 7392 7500 8392 7528
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7429 5963 7463
rect 5905 7423 5963 7429
rect 6365 7463 6423 7469
rect 6365 7429 6377 7463
rect 6411 7460 6423 7463
rect 7006 7460 7012 7472
rect 6411 7432 7012 7460
rect 6411 7429 6423 7432
rect 6365 7423 6423 7429
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2774 7392 2780 7404
rect 2639 7364 2780 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 6086 7352 6092 7404
rect 6144 7352 6150 7404
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7101 7395 7159 7401
rect 7101 7392 7113 7395
rect 6779 7364 7113 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 7101 7361 7113 7364
rect 7147 7361 7159 7395
rect 7101 7355 7159 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7392 7392 7420 7500
rect 8386 7488 8392 7500
rect 8444 7528 8450 7540
rect 8570 7528 8576 7540
rect 8444 7500 8576 7528
rect 8444 7488 8450 7500
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 8662 7488 8668 7540
rect 8720 7488 8726 7540
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 8996 7500 9260 7528
rect 8996 7488 9002 7500
rect 7742 7420 7748 7472
rect 7800 7420 7806 7472
rect 8680 7460 8708 7488
rect 8680 7432 9168 7460
rect 7331 7364 7420 7392
rect 7561 7395 7619 7401
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 2038 7284 2044 7336
rect 2096 7284 2102 7336
rect 3050 7284 3056 7336
rect 3108 7284 3114 7336
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 6196 7324 6224 7355
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 5868 7296 6224 7324
rect 6472 7296 6837 7324
rect 5868 7284 5874 7296
rect 2406 7216 2412 7268
rect 2464 7216 2470 7268
rect 2777 7259 2835 7265
rect 2777 7225 2789 7259
rect 2823 7256 2835 7259
rect 6181 7259 6239 7265
rect 2823 7228 4752 7256
rect 2823 7225 2835 7228
rect 2777 7219 2835 7225
rect 3697 7191 3755 7197
rect 3697 7157 3709 7191
rect 3743 7188 3755 7191
rect 4614 7188 4620 7200
rect 3743 7160 4620 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 4724 7188 4752 7228
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 6472 7256 6500 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6227 7228 6500 7256
rect 7116 7256 7144 7355
rect 7576 7324 7604 7355
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 7760 7392 7788 7420
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7760 7364 7849 7392
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8941 7395 8999 7401
rect 8312 7364 8892 7392
rect 8312 7324 8340 7364
rect 7576 7296 8340 7324
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 7116 7228 7788 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 7760 7200 7788 7228
rect 7834 7216 7840 7268
rect 7892 7216 7898 7268
rect 8294 7216 8300 7268
rect 8352 7216 8358 7268
rect 6362 7188 6368 7200
rect 4724 7160 6368 7188
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 7006 7148 7012 7200
rect 7064 7148 7070 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8496 7188 8524 7287
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 8864 7256 8892 7364
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9030 7392 9036 7404
rect 8987 7364 9036 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9140 7401 9168 7432
rect 9232 7401 9260 7500
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 11940 7500 12572 7528
rect 11940 7488 11946 7500
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9364 7432 9505 7460
rect 9364 7420 9370 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9674 7420 9680 7472
rect 9732 7469 9738 7472
rect 9732 7463 9751 7469
rect 9739 7429 9751 7463
rect 9732 7423 9751 7429
rect 11977 7463 12035 7469
rect 11977 7429 11989 7463
rect 12023 7460 12035 7463
rect 12434 7460 12440 7472
rect 12023 7432 12440 7460
rect 12023 7429 12035 7432
rect 11977 7423 12035 7429
rect 9732 7420 9738 7423
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 12544 7401 12572 7500
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12676 7500 12817 7528
rect 12676 7488 12682 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 15562 7488 15568 7540
rect 15620 7488 15626 7540
rect 16574 7528 16580 7540
rect 15764 7500 16580 7528
rect 14090 7420 14096 7472
rect 14148 7460 14154 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 14148 7432 15025 7460
rect 14148 7420 14154 7432
rect 15013 7429 15025 7432
rect 15059 7460 15071 7463
rect 15764 7460 15792 7500
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 17000 7500 17325 7528
rect 17000 7488 17006 7500
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 17313 7491 17371 7497
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18506 7528 18512 7540
rect 18012 7500 18512 7528
rect 18012 7488 18018 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21048 7500 22416 7528
rect 21048 7488 21054 7500
rect 15059 7432 15792 7460
rect 15841 7463 15899 7469
rect 15059 7429 15071 7432
rect 15013 7423 15071 7429
rect 15841 7429 15853 7463
rect 15887 7460 15899 7463
rect 16206 7460 16212 7472
rect 15887 7432 16212 7460
rect 15887 7429 15899 7432
rect 15841 7423 15899 7429
rect 16206 7420 16212 7432
rect 16264 7460 16270 7472
rect 16264 7432 17448 7460
rect 16264 7420 16270 7432
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 9217 7355 9275 7361
rect 11992 7364 12357 7392
rect 11992 7336 12020 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 15654 7392 15660 7404
rect 12667 7364 15660 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 17420 7401 17448 7432
rect 22186 7420 22192 7472
rect 22244 7420 22250 7472
rect 22278 7420 22284 7472
rect 22336 7420 22342 7472
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18046 7392 18052 7404
rect 18003 7364 18052 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 11974 7284 11980 7336
rect 12032 7284 12038 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 12124 7296 12173 7324
rect 12124 7284 12130 7296
rect 12161 7293 12173 7296
rect 12207 7324 12219 7327
rect 12250 7324 12256 7336
rect 12207 7296 12256 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7324 15531 7327
rect 15764 7324 15792 7355
rect 15519 7296 15792 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 16298 7324 16304 7336
rect 15988 7296 16304 7324
rect 15988 7284 15994 7296
rect 16298 7284 16304 7296
rect 16356 7324 16362 7336
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 16356 7296 16681 7324
rect 16356 7284 16362 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 17972 7324 18000 7355
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 18966 7352 18972 7404
rect 19024 7352 19030 7404
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21407 7364 21864 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 16669 7287 16727 7293
rect 17144 7296 18000 7324
rect 18156 7324 18184 7352
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 18156 7296 18245 7324
rect 9401 7259 9459 7265
rect 9401 7256 9413 7259
rect 8864 7228 9413 7256
rect 9401 7225 9413 7228
rect 9447 7225 9459 7259
rect 9401 7219 9459 7225
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 13446 7256 13452 7268
rect 11940 7228 13452 7256
rect 11940 7216 11946 7228
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 15102 7216 15108 7268
rect 15160 7216 15166 7268
rect 15378 7216 15384 7268
rect 15436 7216 15442 7268
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 17144 7256 17172 7296
rect 18233 7293 18245 7296
rect 18279 7324 18291 7327
rect 18322 7324 18328 7336
rect 18279 7296 18328 7324
rect 18279 7293 18291 7296
rect 18233 7287 18291 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 16163 7228 17172 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 7800 7160 8524 7188
rect 7800 7148 7806 7160
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 8720 7160 8953 7188
rect 8720 7148 8726 7160
rect 8941 7157 8953 7160
rect 8987 7157 8999 7191
rect 8941 7151 8999 7157
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9180 7160 9689 7188
rect 9180 7148 9186 7160
rect 9677 7157 9689 7160
rect 9723 7157 9735 7191
rect 9677 7151 9735 7157
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11606 7188 11612 7200
rect 11563 7160 11612 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 12621 7191 12679 7197
rect 12621 7157 12633 7191
rect 12667 7188 12679 7191
rect 15010 7188 15016 7200
rect 12667 7160 15016 7188
rect 12667 7157 12679 7160
rect 12621 7151 12679 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15120 7188 15148 7216
rect 16132 7188 16160 7219
rect 15120 7160 16160 7188
rect 16298 7148 16304 7200
rect 16356 7148 16362 7200
rect 17144 7188 17172 7228
rect 17402 7216 17408 7268
rect 17460 7256 17466 7268
rect 18141 7259 18199 7265
rect 18141 7256 18153 7259
rect 17460 7228 18153 7256
rect 17460 7216 17466 7228
rect 18141 7225 18153 7228
rect 18187 7225 18199 7259
rect 19904 7256 19932 7352
rect 21836 7265 21864 7364
rect 22388 7333 22416 7500
rect 23106 7420 23112 7472
rect 23164 7460 23170 7472
rect 25133 7463 25191 7469
rect 25133 7460 25145 7463
rect 23164 7432 25145 7460
rect 23164 7420 23170 7432
rect 25133 7429 25145 7432
rect 25179 7429 25191 7463
rect 25133 7423 25191 7429
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 18141 7219 18199 7225
rect 18248 7228 19932 7256
rect 21821 7259 21879 7265
rect 17497 7191 17555 7197
rect 17497 7188 17509 7191
rect 17144 7160 17509 7188
rect 17497 7157 17509 7160
rect 17543 7157 17555 7191
rect 17497 7151 17555 7157
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 17865 7191 17923 7197
rect 17865 7188 17877 7191
rect 17736 7160 17877 7188
rect 17736 7148 17742 7160
rect 17865 7157 17877 7160
rect 17911 7157 17923 7191
rect 17865 7151 17923 7157
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18248 7188 18276 7228
rect 21821 7225 21833 7259
rect 21867 7225 21879 7259
rect 21821 7219 21879 7225
rect 18095 7160 18276 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18322 7148 18328 7200
rect 18380 7148 18386 7200
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19334 7188 19340 7200
rect 18831 7160 19340 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 21174 7148 21180 7200
rect 21232 7148 21238 7200
rect 25409 7191 25467 7197
rect 25409 7157 25421 7191
rect 25455 7188 25467 7191
rect 25455 7160 26004 7188
rect 25455 7157 25467 7160
rect 25409 7151 25467 7157
rect 1104 7098 25852 7120
rect 1104 7046 4043 7098
rect 4095 7046 4107 7098
rect 4159 7046 4171 7098
rect 4223 7046 4235 7098
rect 4287 7046 4299 7098
rect 4351 7046 10230 7098
rect 10282 7046 10294 7098
rect 10346 7046 10358 7098
rect 10410 7046 10422 7098
rect 10474 7046 10486 7098
rect 10538 7046 16417 7098
rect 16469 7046 16481 7098
rect 16533 7046 16545 7098
rect 16597 7046 16609 7098
rect 16661 7046 16673 7098
rect 16725 7046 22604 7098
rect 22656 7046 22668 7098
rect 22720 7046 22732 7098
rect 22784 7046 22796 7098
rect 22848 7046 22860 7098
rect 22912 7046 25852 7098
rect 1104 7024 25852 7046
rect 25976 6996 26004 7160
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7834 6984 7840 6996
rect 7423 6956 7840 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 8662 6984 8668 6996
rect 7944 6956 8668 6984
rect 4157 6919 4215 6925
rect 4157 6885 4169 6919
rect 4203 6885 4215 6919
rect 4157 6879 4215 6885
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 4706 6916 4712 6928
rect 4571 6888 4712 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 4172 6848 4200 6879
rect 4706 6876 4712 6888
rect 4764 6876 4770 6928
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6885 5135 6919
rect 5077 6879 5135 6885
rect 5092 6848 5120 6879
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 6822 6916 6828 6928
rect 6144 6888 6828 6916
rect 6144 6876 6150 6888
rect 6822 6876 6828 6888
rect 6880 6916 6886 6928
rect 7944 6916 7972 6956
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 8846 6944 8852 6996
rect 8904 6984 8910 6996
rect 9122 6984 9128 6996
rect 8904 6956 9128 6984
rect 8904 6944 8910 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 10137 6987 10195 6993
rect 9272 6956 9536 6984
rect 9272 6944 9278 6956
rect 6880 6888 7972 6916
rect 8128 6888 8984 6916
rect 6880 6876 6886 6888
rect 2464 6820 5120 6848
rect 5261 6851 5319 6857
rect 2464 6808 2470 6820
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5307 6820 5764 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 3844 6752 4445 6780
rect 3844 6740 3850 6752
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5350 6780 5356 6792
rect 4663 6752 5356 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6782 5687 6783
rect 5736 6782 5764 6820
rect 6270 6808 6276 6860
rect 6328 6808 6334 6860
rect 5675 6754 5764 6782
rect 5675 6749 5687 6754
rect 5629 6743 5687 6749
rect 2038 6672 2044 6724
rect 2096 6712 2102 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 2096 6684 3893 6712
rect 2096 6672 2102 6684
rect 3881 6681 3893 6684
rect 3927 6712 3939 6715
rect 4801 6715 4859 6721
rect 4801 6712 4813 6715
rect 3927 6684 4813 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4801 6681 4813 6684
rect 4847 6712 4859 6715
rect 6288 6712 6316 6808
rect 6840 6789 6868 6876
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 8128 6848 8156 6888
rect 7699 6820 8156 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8754 6808 8760 6860
rect 8812 6808 8818 6860
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6972 6752 7021 6780
rect 6972 6740 6978 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7098 6740 7104 6792
rect 7156 6740 7162 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7837 6743 7895 6749
rect 7944 6752 8217 6780
rect 4847 6684 6316 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 7466 6672 7472 6724
rect 7524 6712 7530 6724
rect 7852 6712 7880 6743
rect 7524 6684 7880 6712
rect 7524 6672 7530 6684
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 5350 6644 5356 6656
rect 4387 6616 5356 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 7834 6644 7840 6656
rect 6687 6616 7840 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 7834 6604 7840 6616
rect 7892 6644 7898 6656
rect 7944 6644 7972 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 8772 6780 8800 6808
rect 8956 6789 8984 6888
rect 9398 6876 9404 6928
rect 9456 6876 9462 6928
rect 9508 6916 9536 6956
rect 10137 6953 10149 6987
rect 10183 6953 10195 6987
rect 10137 6947 10195 6953
rect 9861 6919 9919 6925
rect 9508 6888 9720 6916
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9692 6848 9720 6888
rect 9861 6885 9873 6919
rect 9907 6916 9919 6919
rect 10152 6916 10180 6947
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12492 6956 13185 6984
rect 12492 6944 12498 6956
rect 13173 6953 13185 6956
rect 13219 6984 13231 6987
rect 14274 6984 14280 6996
rect 13219 6956 14280 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15010 6944 15016 6996
rect 15068 6984 15074 6996
rect 18046 6984 18052 6996
rect 15068 6956 18052 6984
rect 15068 6944 15074 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18233 6987 18291 6993
rect 18233 6953 18245 6987
rect 18279 6984 18291 6987
rect 18506 6984 18512 6996
rect 18279 6956 18512 6984
rect 18279 6953 18291 6956
rect 18233 6947 18291 6953
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 18966 6944 18972 6996
rect 19024 6944 19030 6996
rect 25958 6944 25964 6996
rect 26016 6944 26022 6996
rect 10778 6916 10784 6928
rect 9907 6888 10784 6916
rect 9907 6885 9919 6888
rect 9861 6879 9919 6885
rect 10778 6876 10784 6888
rect 10836 6876 10842 6928
rect 11241 6919 11299 6925
rect 11241 6885 11253 6919
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9539 6820 9628 6848
rect 9692 6820 9965 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 8711 6752 8800 6780
rect 8941 6783 8999 6789
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 8941 6749 8953 6783
rect 8987 6780 8999 6783
rect 9122 6780 9128 6792
rect 8987 6752 9128 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 8496 6712 8524 6740
rect 8352 6684 8524 6712
rect 8588 6712 8616 6743
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9306 6780 9312 6792
rect 9180 6752 9312 6780
rect 9180 6740 9186 6752
rect 9306 6740 9312 6752
rect 9364 6780 9370 6792
rect 9600 6780 9628 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 11256 6848 11284 6879
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 17954 6916 17960 6928
rect 15436 6888 17960 6916
rect 15436 6876 15442 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6916 18199 6919
rect 18984 6916 19012 6944
rect 18187 6888 19012 6916
rect 20257 6919 20315 6925
rect 18187 6885 18199 6888
rect 18141 6879 18199 6885
rect 20257 6885 20269 6919
rect 20303 6885 20315 6919
rect 20257 6879 20315 6885
rect 11330 6848 11336 6860
rect 11256 6820 11336 6848
rect 9953 6811 10011 6817
rect 11330 6808 11336 6820
rect 11388 6848 11394 6860
rect 12066 6848 12072 6860
rect 11388 6820 12072 6848
rect 11388 6808 11394 6820
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 12308 6820 18797 6848
rect 12308 6808 12314 6820
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 19337 6851 19395 6857
rect 19337 6817 19349 6851
rect 19383 6848 19395 6851
rect 19794 6848 19800 6860
rect 19383 6820 19800 6848
rect 19383 6817 19395 6820
rect 19337 6811 19395 6817
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20272 6848 20300 6879
rect 19852 6820 20300 6848
rect 22281 6851 22339 6857
rect 19852 6808 19858 6820
rect 22281 6817 22293 6851
rect 22327 6848 22339 6851
rect 22370 6848 22376 6860
rect 22327 6820 22376 6848
rect 22327 6817 22339 6820
rect 22281 6811 22339 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 9766 6780 9772 6792
rect 9364 6752 9536 6780
rect 9600 6752 9772 6780
rect 9364 6740 9370 6752
rect 9030 6712 9036 6724
rect 8588 6684 9036 6712
rect 8352 6672 8358 6684
rect 9030 6672 9036 6684
rect 9088 6712 9094 6724
rect 9398 6712 9404 6724
rect 9088 6684 9404 6712
rect 9088 6672 9094 6684
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 9508 6712 9536 6752
rect 9766 6740 9772 6752
rect 9824 6780 9830 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9824 6752 10057 6780
rect 9824 6740 9830 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 11238 6740 11244 6792
rect 11296 6780 11302 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11296 6752 11437 6780
rect 11296 6740 11302 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 16577 6783 16635 6789
rect 16577 6780 16589 6783
rect 16264 6752 16589 6780
rect 16264 6740 16270 6752
rect 16577 6749 16589 6752
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 16942 6780 16948 6792
rect 16807 6752 16948 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 17770 6780 17776 6792
rect 17727 6752 17776 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18104 6752 18613 6780
rect 18104 6740 18110 6752
rect 18601 6749 18613 6752
rect 18647 6780 18659 6783
rect 18966 6780 18972 6792
rect 18647 6752 18972 6780
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 20530 6740 20536 6792
rect 20588 6740 20594 6792
rect 10873 6715 10931 6721
rect 9508 6684 10548 6712
rect 7892 6616 7972 6644
rect 8021 6647 8079 6653
rect 7892 6604 7898 6616
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 9674 6644 9680 6656
rect 8067 6616 9680 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10520 6653 10548 6684
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 10919 6684 11652 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 10505 6647 10563 6653
rect 10505 6613 10517 6647
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 11330 6604 11336 6656
rect 11388 6604 11394 6656
rect 11624 6644 11652 6684
rect 11698 6672 11704 6724
rect 11756 6672 11762 6724
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 15654 6672 15660 6724
rect 15712 6712 15718 6724
rect 16298 6712 16304 6724
rect 15712 6684 16304 6712
rect 15712 6672 15718 6684
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 19981 6715 20039 6721
rect 19981 6712 19993 6715
rect 19300 6684 19993 6712
rect 19300 6672 19306 6684
rect 19981 6681 19993 6684
rect 20027 6712 20039 6715
rect 20027 6684 20576 6712
rect 20027 6681 20039 6684
rect 19981 6675 20039 6681
rect 11882 6644 11888 6656
rect 11624 6616 11888 6644
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16945 6647 17003 6653
rect 16945 6644 16957 6647
rect 16172 6616 16957 6644
rect 16172 6604 16178 6616
rect 16945 6613 16957 6616
rect 16991 6613 17003 6647
rect 16945 6607 17003 6613
rect 18693 6647 18751 6653
rect 18693 6613 18705 6647
rect 18739 6644 18751 6647
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 18739 6616 19901 6644
rect 18739 6613 18751 6616
rect 18693 6607 18751 6613
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 20441 6647 20499 6653
rect 20441 6644 20453 6647
rect 20128 6616 20453 6644
rect 20128 6604 20134 6616
rect 20441 6613 20453 6616
rect 20487 6613 20499 6647
rect 20548 6644 20576 6684
rect 20806 6672 20812 6724
rect 20864 6672 20870 6724
rect 21450 6672 21456 6724
rect 21508 6672 21514 6724
rect 20714 6644 20720 6656
rect 20548 6616 20720 6644
rect 20441 6607 20499 6613
rect 20714 6604 20720 6616
rect 20772 6644 20778 6656
rect 21726 6644 21732 6656
rect 20772 6616 21732 6644
rect 20772 6604 20778 6616
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 1104 6554 25852 6576
rect 1104 6502 4703 6554
rect 4755 6502 4767 6554
rect 4819 6502 4831 6554
rect 4883 6502 4895 6554
rect 4947 6502 4959 6554
rect 5011 6502 10890 6554
rect 10942 6502 10954 6554
rect 11006 6502 11018 6554
rect 11070 6502 11082 6554
rect 11134 6502 11146 6554
rect 11198 6502 17077 6554
rect 17129 6502 17141 6554
rect 17193 6502 17205 6554
rect 17257 6502 17269 6554
rect 17321 6502 17333 6554
rect 17385 6502 23264 6554
rect 23316 6502 23328 6554
rect 23380 6502 23392 6554
rect 23444 6502 23456 6554
rect 23508 6502 23520 6554
rect 23572 6502 25852 6554
rect 1104 6480 25852 6502
rect 4632 6412 5764 6440
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 4632 6313 4660 6412
rect 4908 6344 5488 6372
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4706 6264 4712 6316
rect 4764 6264 4770 6316
rect 4908 6313 4936 6344
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6306 5227 6307
rect 5215 6304 5304 6306
rect 5350 6304 5356 6316
rect 5215 6278 5356 6304
rect 5215 6273 5227 6278
rect 5276 6276 5356 6278
rect 5169 6267 5227 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 5460 6236 5488 6344
rect 5736 6316 5764 6412
rect 7006 6400 7012 6452
rect 7064 6400 7070 6452
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7800 6412 7941 6440
rect 7800 6400 7806 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 8754 6440 8760 6452
rect 8496 6412 8760 6440
rect 7024 6372 7052 6400
rect 5828 6344 7052 6372
rect 7208 6372 7236 6400
rect 8205 6375 8263 6381
rect 7208 6344 8156 6372
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 5828 6313 5856 6344
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6178 6304 6184 6316
rect 6043 6276 6184 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 6012 6236 6040 6267
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6564 6276 6837 6304
rect 5460 6208 6040 6236
rect 2700 6168 2728 6196
rect 6564 6168 6592 6276
rect 6825 6273 6837 6276
rect 6871 6304 6883 6307
rect 7006 6304 7012 6316
rect 6871 6276 7012 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 8128 6313 8156 6344
rect 8205 6341 8217 6375
rect 8251 6372 8263 6375
rect 8312 6372 8340 6400
rect 8251 6344 8340 6372
rect 8251 6341 8263 6344
rect 8205 6335 8263 6341
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 7024 6236 7052 6264
rect 7837 6239 7895 6245
rect 7024 6208 7788 6236
rect 2700 6140 6592 6168
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 7331 6140 7696 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 7668 6112 7696 6140
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4614 6100 4620 6112
rect 4295 6072 4620 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 4985 6103 5043 6109
rect 4985 6069 4997 6103
rect 5031 6100 5043 6103
rect 5074 6100 5080 6112
rect 5031 6072 5080 6100
rect 5031 6069 5043 6072
rect 4985 6063 5043 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5258 6060 5264 6112
rect 5316 6100 5322 6112
rect 5353 6103 5411 6109
rect 5353 6100 5365 6103
rect 5316 6072 5365 6100
rect 5316 6060 5322 6072
rect 5353 6069 5365 6072
rect 5399 6069 5411 6103
rect 5353 6063 5411 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6788 6072 6929 6100
rect 6788 6060 6794 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7558 6060 7564 6112
rect 7616 6060 7622 6112
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 7760 6100 7788 6208
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8220 6236 8248 6335
rect 8386 6332 8392 6384
rect 8444 6332 8450 6384
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8404 6304 8432 6332
rect 8496 6313 8524 6412
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11698 6440 11704 6452
rect 11563 6412 11704 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11882 6400 11888 6452
rect 11940 6400 11946 6452
rect 12342 6400 12348 6452
rect 12400 6400 12406 6452
rect 14826 6400 14832 6452
rect 14884 6400 14890 6452
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 15838 6400 15844 6452
rect 15896 6400 15902 6452
rect 16298 6400 16304 6452
rect 16356 6400 16362 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16448 6412 19656 6440
rect 16448 6400 16454 6412
rect 9232 6372 9260 6400
rect 9692 6372 9720 6400
rect 8588 6344 9260 6372
rect 9324 6344 9720 6372
rect 8588 6313 8616 6344
rect 8343 6276 8432 6304
rect 8481 6307 8539 6313
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9324 6304 9352 6344
rect 11606 6332 11612 6384
rect 11664 6332 11670 6384
rect 11793 6375 11851 6381
rect 11793 6341 11805 6375
rect 11839 6372 11851 6375
rect 11900 6372 11928 6400
rect 14090 6372 14096 6384
rect 11839 6344 14096 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 15197 6375 15255 6381
rect 15197 6372 15209 6375
rect 14200 6344 15209 6372
rect 9263 6276 9352 6304
rect 9401 6307 9459 6313
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 7883 6208 8248 6236
rect 8757 6239 8815 6245
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 9416 6236 9444 6267
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 9858 6264 9864 6316
rect 9916 6264 9922 6316
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10686 6304 10692 6316
rect 10284 6276 10692 6304
rect 10284 6264 10290 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 11624 6304 11652 6332
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11624 6276 11713 6304
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 11701 6267 11759 6273
rect 12406 6276 12541 6304
rect 8803 6208 9444 6236
rect 9493 6239 9551 6245
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9539 6208 9965 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6205 10103 6239
rect 10045 6199 10103 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12406 6236 12434 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 14200 6245 14228 6344
rect 15197 6341 15209 6344
rect 15243 6341 15255 6375
rect 15197 6335 15255 6341
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 12299 6208 12434 6236
rect 14185 6239 14243 6245
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10060 6168 10088 6199
rect 9732 6140 10088 6168
rect 9732 6128 9738 6140
rect 12066 6128 12072 6180
rect 12124 6128 12130 6180
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 13906 6168 13912 6180
rect 12216 6140 13912 6168
rect 12216 6128 12222 6140
rect 13906 6128 13912 6140
rect 13964 6168 13970 6180
rect 14200 6168 14228 6199
rect 14384 6180 14412 6267
rect 15028 6236 15056 6267
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15672 6304 15700 6400
rect 15856 6372 15884 6400
rect 16316 6372 16344 6400
rect 16669 6375 16727 6381
rect 16669 6372 16681 6375
rect 15856 6344 15976 6372
rect 16316 6344 16681 6372
rect 15948 6313 15976 6344
rect 16669 6341 16681 6344
rect 16715 6341 16727 6375
rect 16669 6335 16727 6341
rect 18046 6332 18052 6384
rect 18104 6332 18110 6384
rect 18322 6332 18328 6384
rect 18380 6332 18386 6384
rect 19334 6332 19340 6384
rect 19392 6332 19398 6384
rect 19628 6372 19656 6412
rect 19794 6400 19800 6452
rect 19852 6400 19858 6452
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 20806 6440 20812 6452
rect 20671 6412 20812 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21450 6400 21456 6452
rect 21508 6400 21514 6452
rect 19628 6344 21312 6372
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15672 6276 15853 6304
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 15934 6307 15992 6313
rect 15934 6273 15946 6307
rect 15980 6273 15992 6307
rect 15934 6267 15992 6273
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 15028 6208 15700 6236
rect 13964 6140 14228 6168
rect 13964 6128 13970 6140
rect 14366 6128 14372 6180
rect 14424 6128 14430 6180
rect 14476 6140 14964 6168
rect 10226 6100 10232 6112
rect 7760 6072 10232 6100
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 11422 6100 11428 6112
rect 10459 6072 11428 6100
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 14476 6100 14504 6140
rect 13688 6072 14504 6100
rect 14553 6103 14611 6109
rect 13688 6060 13694 6072
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14826 6100 14832 6112
rect 14599 6072 14832 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 14936 6100 14964 6140
rect 15010 6128 15016 6180
rect 15068 6168 15074 6180
rect 15562 6168 15568 6180
rect 15068 6140 15568 6168
rect 15068 6128 15074 6140
rect 15562 6128 15568 6140
rect 15620 6128 15626 6180
rect 15672 6168 15700 6208
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16132 6236 16160 6264
rect 15804 6208 16160 6236
rect 16224 6236 16252 6267
rect 16298 6264 16304 6316
rect 16356 6313 16362 6316
rect 16356 6267 16364 6313
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 18064 6304 18092 6332
rect 17635 6276 18092 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 16356 6264 16362 6267
rect 20346 6264 20352 6316
rect 20404 6264 20410 6316
rect 20806 6264 20812 6316
rect 20864 6264 20870 6316
rect 16224 6208 16620 6236
rect 15804 6196 15810 6208
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 15672 6140 16497 6168
rect 16485 6137 16497 6140
rect 16531 6137 16543 6171
rect 16592 6168 16620 6208
rect 17310 6196 17316 6248
rect 17368 6236 17374 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 17368 6208 17509 6236
rect 17368 6196 17374 6208
rect 17497 6205 17509 6208
rect 17543 6205 17555 6239
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17497 6199 17555 6205
rect 17972 6208 18061 6236
rect 17972 6180 18000 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18414 6236 18420 6248
rect 18049 6199 18107 6205
rect 18156 6208 18420 6236
rect 17037 6171 17095 6177
rect 17037 6168 17049 6171
rect 16592 6140 17049 6168
rect 16485 6131 16543 6137
rect 17037 6137 17049 6140
rect 17083 6168 17095 6171
rect 17678 6168 17684 6180
rect 17083 6140 17684 6168
rect 17083 6137 17095 6140
rect 17037 6131 17095 6137
rect 17678 6128 17684 6140
rect 17736 6128 17742 6180
rect 17954 6128 17960 6180
rect 18012 6128 18018 6180
rect 16390 6100 16396 6112
rect 14936 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17126 6060 17132 6112
rect 17184 6060 17190 6112
rect 17865 6103 17923 6109
rect 17865 6069 17877 6103
rect 17911 6100 17923 6103
rect 18156 6100 18184 6208
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 20364 6236 20392 6264
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 20364 6208 20913 6236
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 20901 6199 20959 6205
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 21177 6171 21235 6177
rect 21177 6168 21189 6171
rect 20496 6140 21189 6168
rect 20496 6128 20502 6140
rect 21177 6137 21189 6140
rect 21223 6137 21235 6171
rect 21284 6168 21312 6344
rect 21637 6307 21695 6313
rect 21637 6304 21649 6307
rect 21376 6276 21649 6304
rect 21376 6245 21404 6276
rect 21637 6273 21649 6276
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 21726 6264 21732 6316
rect 21784 6304 21790 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21784 6276 22017 6304
rect 21784 6264 21790 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6304 25283 6307
rect 25498 6304 25504 6316
rect 25271 6276 25504 6304
rect 25271 6273 25283 6276
rect 25225 6267 25283 6273
rect 25498 6264 25504 6276
rect 25556 6264 25562 6316
rect 21361 6239 21419 6245
rect 21361 6205 21373 6239
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 24118 6168 24124 6180
rect 21284 6140 24124 6168
rect 21177 6131 21235 6137
rect 24118 6128 24124 6140
rect 24176 6128 24182 6180
rect 25406 6128 25412 6180
rect 25464 6128 25470 6180
rect 17911 6072 18184 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 21818 6060 21824 6112
rect 21876 6060 21882 6112
rect 22370 6060 22376 6112
rect 22428 6100 22434 6112
rect 22830 6100 22836 6112
rect 22428 6072 22836 6100
rect 22428 6060 22434 6072
rect 22830 6060 22836 6072
rect 22888 6060 22894 6112
rect 1104 6010 25852 6032
rect 1104 5958 4043 6010
rect 4095 5958 4107 6010
rect 4159 5958 4171 6010
rect 4223 5958 4235 6010
rect 4287 5958 4299 6010
rect 4351 5958 10230 6010
rect 10282 5958 10294 6010
rect 10346 5958 10358 6010
rect 10410 5958 10422 6010
rect 10474 5958 10486 6010
rect 10538 5958 16417 6010
rect 16469 5958 16481 6010
rect 16533 5958 16545 6010
rect 16597 5958 16609 6010
rect 16661 5958 16673 6010
rect 16725 5958 22604 6010
rect 22656 5958 22668 6010
rect 22720 5958 22732 6010
rect 22784 5958 22796 6010
rect 22848 5958 22860 6010
rect 22912 5958 25852 6010
rect 1104 5936 25852 5958
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5896 6699 5899
rect 7374 5896 7380 5908
rect 6687 5868 7380 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 8573 5899 8631 5905
rect 7616 5868 8432 5896
rect 7616 5856 7622 5868
rect 6730 5788 6736 5840
rect 6788 5828 6794 5840
rect 7285 5831 7343 5837
rect 7285 5828 7297 5831
rect 6788 5800 7297 5828
rect 6788 5788 6794 5800
rect 7285 5797 7297 5800
rect 7331 5797 7343 5831
rect 7285 5791 7343 5797
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5760 5227 5763
rect 5258 5760 5264 5772
rect 5215 5732 5264 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 7006 5720 7012 5772
rect 7064 5720 7070 5772
rect 7484 5760 7512 5856
rect 7650 5788 7656 5840
rect 7708 5828 7714 5840
rect 8404 5837 8432 5868
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8754 5896 8760 5908
rect 8619 5868 8760 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 11330 5856 11336 5908
rect 11388 5856 11394 5908
rect 13906 5856 13912 5908
rect 13964 5856 13970 5908
rect 15194 5896 15200 5908
rect 14568 5868 15200 5896
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7708 5800 7849 5828
rect 7708 5788 7714 5800
rect 7837 5797 7849 5800
rect 7883 5797 7895 5831
rect 7837 5791 7895 5797
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 9398 5828 9404 5840
rect 8435 5800 9404 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 7484 5732 7573 5760
rect 7561 5729 7573 5732
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4488 5664 4905 5692
rect 4488 5652 4494 5664
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 11348 5692 11376 5856
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 4893 5655 4951 5661
rect 6932 5664 8248 5692
rect 11348 5664 11805 5692
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 1535 5596 2774 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 2746 5556 2774 5596
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6932 5624 6960 5664
rect 5500 5596 5658 5624
rect 6472 5596 6960 5624
rect 5500 5584 5506 5596
rect 6472 5556 6500 5596
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 7432 5596 8125 5624
rect 7432 5584 7438 5596
rect 8113 5593 8125 5596
rect 8159 5593 8171 5627
rect 8220 5624 8248 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 13924 5701 13952 5856
rect 14568 5837 14596 5868
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 15286 5856 15292 5908
rect 15344 5856 15350 5908
rect 15381 5899 15439 5905
rect 15381 5865 15393 5899
rect 15427 5896 15439 5899
rect 15427 5868 15884 5896
rect 15427 5865 15439 5868
rect 15381 5859 15439 5865
rect 14553 5831 14611 5837
rect 14553 5797 14565 5831
rect 14599 5797 14611 5831
rect 14553 5791 14611 5797
rect 14737 5831 14795 5837
rect 14737 5797 14749 5831
rect 14783 5828 14795 5831
rect 15654 5828 15660 5840
rect 14783 5800 15660 5828
rect 14783 5797 14795 5800
rect 14737 5791 14795 5797
rect 15654 5788 15660 5800
rect 15712 5788 15718 5840
rect 14642 5720 14648 5772
rect 14700 5720 14706 5772
rect 15746 5760 15752 5772
rect 15488 5732 15752 5760
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 14366 5692 14372 5704
rect 13909 5655 13967 5661
rect 14108 5664 14372 5692
rect 13630 5624 13636 5636
rect 8220 5596 13636 5624
rect 8113 5587 8171 5593
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 13740 5624 13768 5652
rect 14108 5624 14136 5664
rect 14366 5652 14372 5664
rect 14424 5692 14430 5704
rect 15488 5702 15516 5732
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 15856 5760 15884 5868
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17218 5896 17224 5908
rect 17000 5868 17224 5896
rect 17000 5856 17006 5868
rect 17218 5856 17224 5868
rect 17276 5896 17282 5908
rect 17865 5899 17923 5905
rect 17865 5896 17877 5899
rect 17276 5868 17877 5896
rect 17276 5856 17282 5868
rect 17865 5865 17877 5868
rect 17911 5865 17923 5899
rect 19794 5896 19800 5908
rect 17865 5859 17923 5865
rect 19260 5868 19800 5896
rect 16853 5831 16911 5837
rect 16853 5828 16865 5831
rect 16408 5800 16865 5828
rect 16408 5769 16436 5800
rect 16853 5797 16865 5800
rect 16899 5797 16911 5831
rect 17126 5828 17132 5840
rect 16853 5791 16911 5797
rect 16960 5800 17132 5828
rect 16393 5763 16451 5769
rect 15856 5732 16160 5760
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14424 5664 14933 5692
rect 14424 5652 14430 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5692 15071 5695
rect 15304 5692 15516 5702
rect 15059 5674 15516 5692
rect 15059 5664 15332 5674
rect 15059 5661 15071 5664
rect 15013 5655 15071 5661
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 13740 5596 14136 5624
rect 14185 5627 14243 5633
rect 14185 5593 14197 5627
rect 14231 5624 14243 5627
rect 14274 5624 14280 5636
rect 14231 5596 14280 5624
rect 14231 5593 14243 5596
rect 14185 5587 14243 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15286 5624 15292 5636
rect 14844 5596 15292 5624
rect 2746 5528 6500 5556
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8938 5556 8944 5568
rect 8067 5528 8944 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 11609 5559 11667 5565
rect 11609 5525 11621 5559
rect 11655 5556 11667 5559
rect 12434 5556 12440 5568
rect 11655 5528 12440 5556
rect 11655 5525 11667 5528
rect 11609 5519 11667 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 13817 5559 13875 5565
rect 13817 5525 13829 5559
rect 13863 5556 13875 5559
rect 14844 5556 14872 5596
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15672 5568 15700 5655
rect 15838 5652 15844 5704
rect 15896 5652 15902 5704
rect 16132 5624 16160 5732
rect 16393 5729 16405 5763
rect 16439 5729 16451 5763
rect 16960 5760 16988 5800
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 19260 5769 19288 5868
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20809 5899 20867 5905
rect 19904 5868 20760 5896
rect 19613 5831 19671 5837
rect 19613 5797 19625 5831
rect 19659 5828 19671 5831
rect 19904 5828 19932 5868
rect 20732 5840 20760 5868
rect 20809 5865 20821 5899
rect 20855 5896 20867 5899
rect 21726 5896 21732 5908
rect 20855 5868 21732 5896
rect 20855 5865 20867 5868
rect 20809 5859 20867 5865
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 19659 5800 19932 5828
rect 19659 5797 19671 5800
rect 19613 5791 19671 5797
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 20625 5831 20683 5837
rect 20625 5828 20637 5831
rect 20496 5800 20637 5828
rect 20496 5788 20502 5800
rect 20625 5797 20637 5800
rect 20671 5797 20683 5831
rect 20625 5791 20683 5797
rect 20714 5788 20720 5840
rect 20772 5788 20778 5840
rect 19245 5763 19303 5769
rect 16393 5723 16451 5729
rect 16776 5732 16988 5760
rect 17144 5732 19012 5760
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16471 5695 16529 5701
rect 16471 5692 16483 5695
rect 16264 5664 16483 5692
rect 16264 5652 16270 5664
rect 16471 5661 16483 5664
rect 16517 5692 16529 5695
rect 16776 5692 16804 5732
rect 17144 5704 17172 5732
rect 16517 5664 16804 5692
rect 17037 5695 17095 5701
rect 16517 5661 16529 5664
rect 16471 5655 16529 5661
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17126 5692 17132 5704
rect 17083 5664 17132 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 17218 5652 17224 5704
rect 17276 5652 17282 5704
rect 17310 5652 17316 5704
rect 17368 5652 17374 5704
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 18046 5692 18052 5704
rect 17819 5664 18052 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 18046 5652 18052 5664
rect 18104 5692 18110 5704
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18104 5664 18889 5692
rect 18104 5652 18110 5664
rect 18877 5661 18889 5664
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 18984 5692 19012 5732
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19245 5723 19303 5729
rect 19352 5732 19717 5760
rect 19352 5692 19380 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 20346 5720 20352 5772
rect 20404 5720 20410 5772
rect 21174 5720 21180 5772
rect 21232 5720 21238 5772
rect 18984 5664 19380 5692
rect 17328 5624 17356 5652
rect 16132 5596 17356 5624
rect 18509 5627 18567 5633
rect 18509 5593 18521 5627
rect 18555 5593 18567 5627
rect 18509 5587 18567 5593
rect 18693 5627 18751 5633
rect 18693 5593 18705 5627
rect 18739 5624 18751 5627
rect 18984 5624 19012 5664
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 20530 5692 20536 5704
rect 19576 5664 20536 5692
rect 19576 5652 19582 5664
rect 20530 5652 20536 5664
rect 20588 5692 20594 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20588 5664 20913 5692
rect 20588 5652 20594 5664
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 20070 5624 20076 5636
rect 18739 5596 19012 5624
rect 19536 5596 20076 5624
rect 18739 5593 18751 5596
rect 18693 5587 18751 5593
rect 13863 5528 14872 5556
rect 15105 5559 15163 5565
rect 13863 5525 13875 5528
rect 13817 5519 13875 5525
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15654 5556 15660 5568
rect 15151 5528 15660 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 16761 5559 16819 5565
rect 16761 5556 16773 5559
rect 16540 5528 16773 5556
rect 16540 5516 16546 5528
rect 16761 5525 16773 5528
rect 16807 5525 16819 5559
rect 18524 5556 18552 5587
rect 19536 5556 19564 5596
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 21818 5584 21824 5636
rect 21876 5584 21882 5636
rect 18524 5528 19564 5556
rect 22649 5559 22707 5565
rect 16761 5519 16819 5525
rect 22649 5525 22661 5559
rect 22695 5556 22707 5559
rect 23106 5556 23112 5568
rect 22695 5528 23112 5556
rect 22695 5525 22707 5528
rect 22649 5519 22707 5525
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 1104 5466 25852 5488
rect 1104 5414 4703 5466
rect 4755 5414 4767 5466
rect 4819 5414 4831 5466
rect 4883 5414 4895 5466
rect 4947 5414 4959 5466
rect 5011 5414 10890 5466
rect 10942 5414 10954 5466
rect 11006 5414 11018 5466
rect 11070 5414 11082 5466
rect 11134 5414 11146 5466
rect 11198 5414 17077 5466
rect 17129 5414 17141 5466
rect 17193 5414 17205 5466
rect 17257 5414 17269 5466
rect 17321 5414 17333 5466
rect 17385 5414 23264 5466
rect 23316 5414 23328 5466
rect 23380 5414 23392 5466
rect 23444 5414 23456 5466
rect 23508 5414 23520 5466
rect 23572 5414 25852 5466
rect 1104 5392 25852 5414
rect 4430 5312 4436 5364
rect 4488 5312 4494 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5132 5324 5396 5352
rect 5132 5312 5138 5324
rect 4448 5284 4476 5312
rect 3988 5256 4476 5284
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 3988 5225 4016 5256
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 5368 5202 5396 5324
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 7653 5355 7711 5361
rect 7653 5352 7665 5355
rect 6880 5324 7665 5352
rect 6880 5312 6886 5324
rect 7653 5321 7665 5324
rect 7699 5321 7711 5355
rect 7926 5352 7932 5364
rect 7653 5315 7711 5321
rect 7760 5324 7932 5352
rect 7561 5219 7619 5225
rect 3973 5179 4031 5185
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7650 5216 7656 5228
rect 7607 5188 7656 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 7760 5225 7788 5324
rect 7926 5312 7932 5324
rect 7984 5352 7990 5364
rect 8386 5352 8392 5364
rect 7984 5324 8392 5352
rect 7984 5312 7990 5324
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5321 11207 5355
rect 13998 5352 14004 5364
rect 11149 5315 11207 5321
rect 13924 5324 14004 5352
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 9490 5284 9496 5296
rect 7883 5256 9496 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 11164 5284 11192 5315
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 11164 5256 11805 5284
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 12434 5244 12440 5296
rect 12492 5244 12498 5296
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 11330 5176 11336 5228
rect 11388 5176 11394 5228
rect 13814 5176 13820 5228
rect 13872 5176 13878 5228
rect 13924 5225 13952 5324
rect 13998 5312 14004 5324
rect 14056 5352 14062 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 14056 5324 16405 5352
rect 14056 5312 14062 5324
rect 15381 5287 15439 5293
rect 15381 5284 15393 5287
rect 14016 5256 15393 5284
rect 14016 5225 14044 5256
rect 15381 5253 15393 5256
rect 15427 5253 15439 5287
rect 15381 5247 15439 5253
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5216 14243 5219
rect 14458 5216 14464 5228
rect 14231 5188 14464 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4614 5148 4620 5160
rect 4295 5120 4620 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11296 5120 11529 5148
rect 11296 5108 11302 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 14660 5080 14688 5179
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14884 5188 15117 5216
rect 14884 5176 14890 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15286 5216 15292 5228
rect 15243 5188 15292 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15470 5182 15476 5234
rect 15528 5216 15534 5234
rect 15856 5225 15884 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 16942 5352 16948 5364
rect 16816 5324 16948 5352
rect 16816 5312 16822 5324
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17862 5312 17868 5364
rect 17920 5352 17926 5364
rect 19518 5352 19524 5364
rect 17920 5324 19524 5352
rect 17920 5312 17926 5324
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20806 5352 20812 5364
rect 20763 5324 20812 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 20916 5324 25268 5352
rect 16209 5287 16267 5293
rect 16209 5253 16221 5287
rect 16255 5284 16267 5287
rect 17402 5284 17408 5296
rect 16255 5256 17408 5284
rect 16255 5253 16267 5256
rect 16209 5247 16267 5253
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 18230 5244 18236 5296
rect 18288 5244 18294 5296
rect 20165 5287 20223 5293
rect 20165 5253 20177 5287
rect 20211 5284 20223 5287
rect 20346 5284 20352 5296
rect 20211 5256 20352 5284
rect 20211 5253 20223 5256
rect 20165 5247 20223 5253
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 15528 5188 15761 5216
rect 15528 5182 15534 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 15381 5151 15439 5157
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 15562 5148 15568 5160
rect 15427 5120 15568 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15948 5148 15976 5179
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 16080 5188 16129 5216
rect 16080 5176 16086 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16482 5176 16488 5228
rect 16540 5176 16546 5228
rect 18782 5176 18788 5228
rect 18840 5216 18846 5228
rect 20916 5216 20944 5324
rect 21821 5287 21879 5293
rect 21821 5284 21833 5287
rect 18840 5188 20944 5216
rect 21008 5256 21833 5284
rect 18840 5176 18846 5188
rect 15948 5120 16344 5148
rect 5276 5052 8064 5080
rect 14660 5052 16068 5080
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 5276 5012 5304 5052
rect 8036 5024 8064 5052
rect 16040 5024 16068 5052
rect 16316 5024 16344 5120
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 21008 5148 21036 5256
rect 21821 5253 21833 5256
rect 21867 5253 21879 5287
rect 21821 5247 21879 5253
rect 21082 5176 21088 5228
rect 21140 5176 21146 5228
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 22094 5216 22100 5228
rect 21223 5188 22100 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 22094 5176 22100 5188
rect 22152 5216 22158 5228
rect 23014 5216 23020 5228
rect 22152 5188 23020 5216
rect 22152 5176 22158 5188
rect 23014 5176 23020 5188
rect 23072 5176 23078 5228
rect 25240 5225 25268 5324
rect 25225 5219 25283 5225
rect 25225 5185 25237 5219
rect 25271 5185 25283 5219
rect 25225 5179 25283 5185
rect 20404 5120 21036 5148
rect 20404 5108 20410 5120
rect 21358 5108 21364 5160
rect 21416 5148 21422 5160
rect 21726 5148 21732 5160
rect 21416 5120 21732 5148
rect 21416 5108 21422 5120
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 20438 5040 20444 5092
rect 20496 5080 20502 5092
rect 22097 5083 22155 5089
rect 22097 5080 22109 5083
rect 20496 5052 22109 5080
rect 20496 5040 20502 5052
rect 22097 5049 22109 5052
rect 22143 5049 22155 5083
rect 22097 5043 22155 5049
rect 1627 4984 5304 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 8018 4972 8024 5024
rect 8076 4972 8082 5024
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 9088 4984 9137 5012
rect 9088 4972 9094 4984
rect 9125 4981 9137 4984
rect 9171 4981 9183 5015
rect 9125 4975 9183 4981
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 5012 13599 5015
rect 14090 5012 14096 5024
rect 13587 4984 14096 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14918 4972 14924 5024
rect 14976 4972 14982 5024
rect 15470 4972 15476 5024
rect 15528 4972 15534 5024
rect 16022 4972 16028 5024
rect 16080 4972 16086 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 16172 4984 16221 5012
rect 16172 4972 16178 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 20622 4972 20628 5024
rect 20680 4972 20686 5024
rect 22278 4972 22284 5024
rect 22336 4972 22342 5024
rect 25406 4972 25412 5024
rect 25464 4972 25470 5024
rect 1104 4922 25852 4944
rect 1104 4870 4043 4922
rect 4095 4870 4107 4922
rect 4159 4870 4171 4922
rect 4223 4870 4235 4922
rect 4287 4870 4299 4922
rect 4351 4870 10230 4922
rect 10282 4870 10294 4922
rect 10346 4870 10358 4922
rect 10410 4870 10422 4922
rect 10474 4870 10486 4922
rect 10538 4870 16417 4922
rect 16469 4870 16481 4922
rect 16533 4870 16545 4922
rect 16597 4870 16609 4922
rect 16661 4870 16673 4922
rect 16725 4870 22604 4922
rect 22656 4870 22668 4922
rect 22720 4870 22732 4922
rect 22784 4870 22796 4922
rect 22848 4870 22860 4922
rect 22912 4870 25852 4922
rect 1104 4848 25852 4870
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4777 7619 4811
rect 7561 4771 7619 4777
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 5776 4576 7481 4604
rect 5776 4564 5782 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7576 4604 7604 4771
rect 7650 4768 7656 4820
rect 7708 4768 7714 4820
rect 7926 4768 7932 4820
rect 7984 4768 7990 4820
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 11241 4811 11299 4817
rect 8435 4780 11192 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 7668 4740 7696 4768
rect 8573 4743 8631 4749
rect 8573 4740 8585 4743
rect 7668 4712 8585 4740
rect 8573 4709 8585 4712
rect 8619 4709 8631 4743
rect 8573 4703 8631 4709
rect 8018 4604 8024 4616
rect 7576 4576 8024 4604
rect 7469 4567 7527 4573
rect 7484 4536 7512 4567
rect 8018 4564 8024 4576
rect 8076 4604 8082 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 8076 4576 8125 4604
rect 8076 4564 8082 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8680 4536 8708 4780
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9784 4712 9873 4740
rect 9784 4616 9812 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 11164 4740 11192 4780
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 11330 4808 11336 4820
rect 11287 4780 11336 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14737 4811 14795 4817
rect 14737 4808 14749 4811
rect 13872 4780 14749 4808
rect 13872 4768 13878 4780
rect 14737 4777 14749 4780
rect 14783 4777 14795 4811
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 14737 4771 14795 4777
rect 14844 4780 15485 4808
rect 12158 4740 12164 4752
rect 11164 4712 12164 4740
rect 9861 4703 9919 4709
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 13541 4743 13599 4749
rect 13541 4740 13553 4743
rect 12768 4712 13553 4740
rect 12768 4700 12774 4712
rect 13541 4709 13553 4712
rect 13587 4709 13599 4743
rect 13541 4703 13599 4709
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10091 4644 10364 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 10336 4613 10364 4644
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 10744 4644 11897 4672
rect 10744 4632 10750 4644
rect 11885 4641 11897 4644
rect 11931 4672 11943 4675
rect 12250 4672 12256 4684
rect 11931 4644 12256 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12894 4672 12900 4684
rect 12667 4644 12900 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12894 4632 12900 4644
rect 12952 4672 12958 4684
rect 13262 4672 13268 4684
rect 12952 4644 13268 4672
rect 12952 4632 12958 4644
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13556 4672 13584 4703
rect 14274 4700 14280 4752
rect 14332 4740 14338 4752
rect 14844 4740 14872 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 15473 4771 15531 4777
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15804 4780 15853 4808
rect 15804 4768 15810 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 16022 4768 16028 4820
rect 16080 4768 16086 4820
rect 16298 4768 16304 4820
rect 16356 4768 16362 4820
rect 18693 4811 18751 4817
rect 18693 4777 18705 4811
rect 18739 4808 18751 4811
rect 19242 4808 19248 4820
rect 18739 4780 19248 4808
rect 18739 4777 18751 4780
rect 18693 4771 18751 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 20622 4768 20628 4820
rect 20680 4768 20686 4820
rect 14332 4712 14872 4740
rect 14332 4700 14338 4712
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 14976 4712 16252 4740
rect 14976 4700 14982 4712
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13556 4644 14105 4672
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14642 4632 14648 4684
rect 14700 4632 14706 4684
rect 14936 4644 15700 4672
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 11974 4604 11980 4616
rect 11655 4576 11980 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 7484 4508 8708 4536
rect 9585 4539 9643 4545
rect 9585 4505 9597 4539
rect 9631 4505 9643 4539
rect 14660 4536 14688 4632
rect 14936 4598 14964 4644
rect 15672 4616 15700 4644
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15804 4644 16160 4672
rect 15804 4632 15810 4644
rect 15013 4607 15071 4613
rect 15013 4598 15025 4607
rect 14936 4573 15025 4598
rect 15059 4573 15071 4607
rect 14936 4570 15071 4573
rect 15013 4567 15071 4570
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4573 15255 4607
rect 15197 4567 15255 4573
rect 15212 4536 15240 4567
rect 15286 4564 15292 4616
rect 15344 4564 15350 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15562 4604 15568 4616
rect 15436 4576 15568 4604
rect 15436 4564 15442 4576
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 16132 4613 16160 4644
rect 16224 4613 16252 4712
rect 16390 4700 16396 4752
rect 16448 4700 16454 4752
rect 16408 4613 16436 4700
rect 17862 4672 17868 4684
rect 16960 4644 17868 4672
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15712 4576 15945 4604
rect 15712 4564 15718 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4573 16267 4607
rect 16209 4567 16267 4573
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16758 4564 16764 4616
rect 16816 4604 16822 4616
rect 16960 4613 16988 4644
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16816 4576 16957 4604
rect 16816 4564 16822 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 20640 4604 20668 4768
rect 21177 4607 21235 4613
rect 21177 4604 21189 4607
rect 20640 4576 21189 4604
rect 16945 4567 17003 4573
rect 21177 4573 21189 4576
rect 21223 4573 21235 4607
rect 21177 4567 21235 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 23106 4604 23112 4616
rect 22051 4576 23112 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 25222 4564 25228 4616
rect 25280 4564 25286 4616
rect 14660 4508 15240 4536
rect 9585 4499 9643 4505
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 9600 4468 9628 4499
rect 15470 4496 15476 4548
rect 15528 4536 15534 4548
rect 17221 4539 17279 4545
rect 17221 4536 17233 4539
rect 15528 4508 17233 4536
rect 15528 4496 15534 4508
rect 17221 4505 17233 4508
rect 17267 4505 17279 4539
rect 17221 4499 17279 4505
rect 17954 4496 17960 4548
rect 18012 4496 18018 4548
rect 7616 4440 9628 4468
rect 10137 4471 10195 4477
rect 7616 4428 7622 4440
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 10318 4468 10324 4480
rect 10183 4440 10324 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 11747 4440 13185 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 13173 4431 13231 4437
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 13906 4468 13912 4480
rect 13771 4440 13912 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 15838 4468 15844 4480
rect 14875 4440 15844 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 20898 4428 20904 4480
rect 20956 4468 20962 4480
rect 20993 4471 21051 4477
rect 20993 4468 21005 4471
rect 20956 4440 21005 4468
rect 20956 4428 20962 4440
rect 20993 4437 21005 4440
rect 21039 4437 21051 4471
rect 20993 4431 21051 4437
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22649 4471 22707 4477
rect 22649 4468 22661 4471
rect 22152 4440 22661 4468
rect 22152 4428 22158 4440
rect 22649 4437 22661 4440
rect 22695 4437 22707 4471
rect 22649 4431 22707 4437
rect 25406 4428 25412 4480
rect 25464 4428 25470 4480
rect 1104 4378 25852 4400
rect 1104 4326 4703 4378
rect 4755 4326 4767 4378
rect 4819 4326 4831 4378
rect 4883 4326 4895 4378
rect 4947 4326 4959 4378
rect 5011 4326 10890 4378
rect 10942 4326 10954 4378
rect 11006 4326 11018 4378
rect 11070 4326 11082 4378
rect 11134 4326 11146 4378
rect 11198 4326 17077 4378
rect 17129 4326 17141 4378
rect 17193 4326 17205 4378
rect 17257 4326 17269 4378
rect 17321 4326 17333 4378
rect 17385 4326 23264 4378
rect 23316 4326 23328 4378
rect 23380 4326 23392 4378
rect 23444 4326 23456 4378
rect 23508 4326 23520 4378
rect 23572 4326 25852 4378
rect 1104 4304 25852 4326
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 11974 4264 11980 4276
rect 5500 4236 11980 4264
rect 5500 4224 5506 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 14274 4224 14280 4276
rect 14332 4224 14338 4276
rect 14734 4224 14740 4276
rect 14792 4224 14798 4276
rect 14826 4224 14832 4276
rect 14884 4224 14890 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 17954 4264 17960 4276
rect 17911 4236 17960 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 22278 4224 22284 4276
rect 22336 4224 22342 4276
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 9582 4196 9588 4208
rect 7984 4168 9588 4196
rect 7984 4156 7990 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 10318 4156 10324 4208
rect 10376 4156 10382 4208
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5592 4100 6377 4128
rect 5592 4088 5598 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4128 7251 4131
rect 7374 4128 7380 4140
rect 7239 4100 7380 4128
rect 7239 4097 7251 4100
rect 7193 4091 7251 4097
rect 5994 4060 6000 4072
rect 5920 4032 6000 4060
rect 5920 4001 5948 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6380 4060 6408 4091
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7515 4100 7788 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7558 4060 7564 4072
rect 6380 4032 7564 4060
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 7760 4060 7788 4100
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8018 4128 8024 4140
rect 7892 4100 8024 4128
rect 7892 4088 7898 4100
rect 8018 4088 8024 4100
rect 8076 4128 8082 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 8076 4100 8125 4128
rect 8076 4088 8082 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 11054 4088 11060 4140
rect 11112 4088 11118 4140
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 8202 4060 8208 4072
rect 7760 4032 8208 4060
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 9030 4060 9036 4072
rect 8352 4032 9036 4060
rect 8352 4020 8358 4032
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 12529 4063 12587 4069
rect 9355 4032 10916 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 6641 3995 6699 4001
rect 6641 3992 6653 3995
rect 5951 3964 6653 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 6641 3961 6653 3964
rect 6687 3992 6699 3995
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 6687 3964 7849 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7837 3961 7849 3964
rect 7883 3992 7895 3995
rect 7926 3992 7932 4004
rect 7883 3964 7932 3992
rect 7883 3961 7895 3964
rect 7837 3955 7895 3961
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 8938 3992 8944 4004
rect 8036 3964 8944 3992
rect 5994 3884 6000 3936
rect 6052 3884 6058 3936
rect 6822 3884 6828 3936
rect 6880 3884 6886 3936
rect 7006 3884 7012 3936
rect 7064 3884 7070 3936
rect 7282 3884 7288 3936
rect 7340 3884 7346 3936
rect 8036 3933 8064 3964
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 10778 3952 10784 4004
rect 10836 3952 10842 4004
rect 10888 4001 10916 4032
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12710 4060 12716 4072
rect 12575 4032 12716 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13740 4060 13768 4091
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14292 4128 14320 4224
rect 14844 4196 14872 4224
rect 14660 4168 14872 4196
rect 14660 4137 14688 4168
rect 20898 4156 20904 4208
rect 20956 4156 20962 4208
rect 14139 4100 14320 4128
rect 14645 4131 14703 4137
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4128 14887 4131
rect 15286 4128 15292 4140
rect 14875 4100 15292 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 13035 4032 13768 4060
rect 13924 4060 13952 4088
rect 14844 4060 14872 4091
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17678 4128 17684 4140
rect 17359 4100 17684 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 13924 4032 14872 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 17328 4060 17356 4091
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 15068 4032 17356 4060
rect 17773 4063 17831 4069
rect 15068 4020 15074 4032
rect 17773 4029 17785 4063
rect 17819 4060 17831 4063
rect 18064 4060 18092 4091
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19576 4100 19901 4128
rect 19576 4088 19582 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22296 4137 22324 4224
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4097 22339 4131
rect 22281 4091 22339 4097
rect 17819 4032 18092 4060
rect 17819 4029 17831 4032
rect 17773 4023 17831 4029
rect 19702 4020 19708 4072
rect 19760 4020 19766 4072
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20211 4032 21864 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 10873 3995 10931 4001
rect 10873 3961 10885 3995
rect 10919 3961 10931 3995
rect 10873 3955 10931 3961
rect 12894 3952 12900 4004
rect 12952 3952 12958 4004
rect 13722 3952 13728 4004
rect 13780 3952 13786 4004
rect 14553 3995 14611 4001
rect 14553 3961 14565 3995
rect 14599 3992 14611 3995
rect 15654 3992 15660 4004
rect 14599 3964 15660 3992
rect 14599 3961 14611 3964
rect 14553 3955 14611 3961
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 17494 3952 17500 4004
rect 17552 3992 17558 4004
rect 17589 3995 17647 4001
rect 17589 3992 17601 3995
rect 17552 3964 17601 3992
rect 17552 3952 17558 3964
rect 17589 3961 17601 3964
rect 17635 3961 17647 3995
rect 17589 3955 17647 3961
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8444 3896 8769 3924
rect 8444 3884 8450 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 10796 3924 10824 3952
rect 9916 3896 10824 3924
rect 9916 3884 9922 3896
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 14185 3927 14243 3933
rect 14185 3924 14197 3927
rect 12676 3896 14197 3924
rect 12676 3884 12682 3896
rect 14185 3893 14197 3896
rect 14231 3924 14243 3927
rect 14274 3924 14280 3936
rect 14231 3896 14280 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 19720 3924 19748 4020
rect 21836 4001 21864 4032
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3961 21879 3995
rect 21821 3955 21879 3961
rect 21637 3927 21695 3933
rect 21637 3924 21649 3927
rect 19720 3896 21649 3924
rect 21637 3893 21649 3896
rect 21683 3893 21695 3927
rect 21637 3887 21695 3893
rect 22097 3927 22155 3933
rect 22097 3893 22109 3927
rect 22143 3924 22155 3927
rect 22278 3924 22284 3936
rect 22143 3896 22284 3924
rect 22143 3893 22155 3896
rect 22097 3887 22155 3893
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 24946 3924 24952 3936
rect 23716 3896 24952 3924
rect 23716 3884 23722 3896
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 1104 3834 25852 3856
rect 1104 3782 4043 3834
rect 4095 3782 4107 3834
rect 4159 3782 4171 3834
rect 4223 3782 4235 3834
rect 4287 3782 4299 3834
rect 4351 3782 10230 3834
rect 10282 3782 10294 3834
rect 10346 3782 10358 3834
rect 10410 3782 10422 3834
rect 10474 3782 10486 3834
rect 10538 3782 16417 3834
rect 16469 3782 16481 3834
rect 16533 3782 16545 3834
rect 16597 3782 16609 3834
rect 16661 3782 16673 3834
rect 16725 3782 22604 3834
rect 22656 3782 22668 3834
rect 22720 3782 22732 3834
rect 22784 3782 22796 3834
rect 22848 3782 22860 3834
rect 22912 3782 25852 3834
rect 1104 3760 25852 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 5258 3720 5264 3732
rect 2179 3692 5264 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6352 3723 6410 3729
rect 6352 3689 6364 3723
rect 6398 3720 6410 3723
rect 7006 3720 7012 3732
rect 6398 3692 7012 3720
rect 6398 3689 6410 3692
rect 6352 3683 6410 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7432 3692 7941 3720
rect 7432 3680 7438 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8260 3692 8953 3720
rect 8260 3680 8266 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 11054 3720 11060 3732
rect 9815 3692 11060 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11228 3723 11286 3729
rect 11228 3689 11240 3723
rect 11274 3720 11286 3723
rect 11422 3720 11428 3732
rect 11274 3692 11428 3720
rect 11274 3689 11286 3692
rect 11228 3683 11286 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 23658 3720 23664 3732
rect 12636 3692 23664 3720
rect 7834 3612 7840 3664
rect 7892 3612 7898 3664
rect 8312 3624 11008 3652
rect 8312 3596 8340 3624
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 4264 3556 6101 3584
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 4264 3525 4292 3556
rect 6089 3553 6101 3556
rect 6135 3584 6147 3587
rect 8294 3584 8300 3596
rect 6135 3556 8300 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8386 3544 8392 3596
rect 8444 3544 8450 3596
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3584 8631 3587
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 8619 3556 9597 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 9585 3553 9597 3556
rect 9631 3584 9643 3587
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 9631 3556 10425 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 10413 3553 10425 3556
rect 10459 3584 10471 3587
rect 10686 3584 10692 3596
rect 10459 3556 10692 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1084 3488 1961 3516
rect 1084 3476 1090 3488
rect 1949 3485 1961 3488
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 1489 3451 1547 3457
rect 1489 3417 1501 3451
rect 1535 3448 1547 3451
rect 4264 3448 4292 3479
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8588 3516 8616 3547
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10980 3593 11008 3624
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11238 3584 11244 3596
rect 11011 3556 11244 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 7800 3488 8616 3516
rect 10137 3519 10195 3525
rect 7800 3476 7806 3488
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10183 3488 10364 3516
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 4430 3448 4436 3460
rect 1535 3420 2774 3448
rect 4264 3420 4436 3448
rect 1535 3417 1547 3420
rect 1489 3411 1547 3417
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 2746 3380 2774 3420
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 4522 3408 4528 3460
rect 4580 3408 4586 3460
rect 4614 3408 4620 3460
rect 4672 3408 4678 3460
rect 5810 3448 5816 3460
rect 5750 3420 5816 3448
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 7098 3408 7104 3460
rect 7156 3408 7162 3460
rect 8297 3451 8355 3457
rect 8297 3417 8309 3451
rect 8343 3448 8355 3451
rect 9122 3448 9128 3460
rect 8343 3420 9128 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 9122 3408 9128 3420
rect 9180 3448 9186 3460
rect 9582 3448 9588 3460
rect 9180 3420 9588 3448
rect 9180 3408 9186 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 10229 3451 10287 3457
rect 10229 3448 10241 3451
rect 9916 3420 10241 3448
rect 9916 3408 9922 3420
rect 10229 3417 10241 3420
rect 10275 3417 10287 3451
rect 10336 3448 10364 3488
rect 10502 3476 10508 3528
rect 10560 3516 10566 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 10560 3488 10793 3516
rect 10560 3476 10566 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 12526 3448 12532 3460
rect 10336 3420 11376 3448
rect 12466 3420 12532 3448
rect 10229 3411 10287 3417
rect 4632 3380 4660 3408
rect 11348 3392 11376 3420
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 2746 3352 4660 3380
rect 5997 3383 6055 3389
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 6730 3380 6736 3392
rect 6043 3352 6736 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3340 9462 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 9824 3352 10609 3380
rect 9824 3340 9830 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 10597 3343 10655 3349
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 12636 3380 12664 3692
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 24762 3680 24768 3732
rect 24820 3680 24826 3732
rect 24854 3680 24860 3732
rect 24912 3720 24918 3732
rect 25041 3723 25099 3729
rect 25041 3720 25053 3723
rect 24912 3692 25053 3720
rect 24912 3680 24918 3692
rect 25041 3689 25053 3692
rect 25087 3689 25099 3723
rect 25041 3683 25099 3689
rect 13173 3655 13231 3661
rect 13173 3621 13185 3655
rect 13219 3652 13231 3655
rect 13354 3652 13360 3664
rect 13219 3624 13360 3652
rect 13219 3621 13231 3624
rect 13173 3615 13231 3621
rect 13354 3612 13360 3624
rect 13412 3652 13418 3664
rect 13630 3652 13636 3664
rect 13412 3624 13636 3652
rect 13412 3612 13418 3624
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 15654 3652 15660 3664
rect 14240 3624 15660 3652
rect 14240 3612 14246 3624
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 24780 3652 24808 3680
rect 25317 3655 25375 3661
rect 25317 3652 25329 3655
rect 24780 3624 25329 3652
rect 25317 3621 25329 3624
rect 25363 3621 25375 3655
rect 25317 3615 25375 3621
rect 15010 3544 15016 3596
rect 15068 3544 15074 3596
rect 16758 3584 16764 3596
rect 15764 3556 16764 3584
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3516 12863 3519
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 12851 3488 13369 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 13357 3485 13369 3488
rect 13403 3516 13415 3519
rect 14550 3516 14556 3528
rect 13403 3488 14556 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 14550 3476 14556 3488
rect 14608 3516 14614 3528
rect 15028 3516 15056 3544
rect 14608 3488 15056 3516
rect 14608 3476 14614 3488
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 15764 3525 15792 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 19576 3556 21005 3584
rect 19576 3544 19582 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 22925 3587 22983 3593
rect 22925 3584 22937 3587
rect 22787 3556 22937 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 22925 3553 22937 3556
rect 22971 3584 22983 3587
rect 24854 3584 24860 3596
rect 22971 3556 24860 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 15764 3448 15792 3479
rect 17770 3476 17776 3528
rect 17828 3476 17834 3528
rect 20898 3476 20904 3528
rect 20956 3476 20962 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22336 3488 22402 3516
rect 22336 3476 22342 3488
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 24670 3516 24676 3528
rect 23072 3488 24676 3516
rect 23072 3476 23078 3488
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 24946 3516 24952 3528
rect 24811 3488 24952 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 25225 3519 25283 3525
rect 25225 3485 25237 3519
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 25958 3516 25964 3528
rect 25547 3488 25964 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 13924 3420 15792 3448
rect 16025 3451 16083 3457
rect 13924 3392 13952 3420
rect 16025 3417 16037 3451
rect 16071 3448 16083 3451
rect 16114 3448 16120 3460
rect 16071 3420 16120 3448
rect 16071 3417 16083 3420
rect 16025 3411 16083 3417
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 17402 3448 17408 3460
rect 17250 3420 17408 3448
rect 17402 3408 17408 3420
rect 17460 3408 17466 3460
rect 21269 3451 21327 3457
rect 21269 3417 21281 3451
rect 21315 3417 21327 3451
rect 25240 3448 25268 3479
rect 25958 3476 25964 3488
rect 26016 3476 26022 3528
rect 25866 3448 25872 3460
rect 21269 3411 21327 3417
rect 22664 3420 24992 3448
rect 25240 3420 25872 3448
rect 11388 3352 12664 3380
rect 11388 3340 11394 3352
rect 12710 3340 12716 3392
rect 12768 3340 12774 3392
rect 13262 3340 13268 3392
rect 13320 3340 13326 3392
rect 13814 3340 13820 3392
rect 13872 3340 13878 3392
rect 13906 3340 13912 3392
rect 13964 3340 13970 3392
rect 14918 3340 14924 3392
rect 14976 3340 14982 3392
rect 20717 3383 20775 3389
rect 20717 3349 20729 3383
rect 20763 3380 20775 3383
rect 21284 3380 21312 3411
rect 20763 3352 21312 3380
rect 20763 3349 20775 3352
rect 20717 3343 20775 3349
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 22664 3380 22692 3420
rect 21600 3352 22692 3380
rect 21600 3340 21606 3352
rect 22830 3340 22836 3392
rect 22888 3380 22894 3392
rect 24964 3389 24992 3420
rect 25866 3408 25872 3420
rect 25924 3408 25930 3460
rect 23477 3383 23535 3389
rect 23477 3380 23489 3383
rect 22888 3352 23489 3380
rect 22888 3340 22894 3352
rect 23477 3349 23489 3352
rect 23523 3349 23535 3383
rect 23477 3343 23535 3349
rect 24949 3383 25007 3389
rect 24949 3349 24961 3383
rect 24995 3349 25007 3383
rect 24949 3343 25007 3349
rect 1104 3290 25852 3312
rect 1104 3238 4703 3290
rect 4755 3238 4767 3290
rect 4819 3238 4831 3290
rect 4883 3238 4895 3290
rect 4947 3238 4959 3290
rect 5011 3238 10890 3290
rect 10942 3238 10954 3290
rect 11006 3238 11018 3290
rect 11070 3238 11082 3290
rect 11134 3238 11146 3290
rect 11198 3238 17077 3290
rect 17129 3238 17141 3290
rect 17193 3238 17205 3290
rect 17257 3238 17269 3290
rect 17321 3238 17333 3290
rect 17385 3238 23264 3290
rect 23316 3238 23328 3290
rect 23380 3238 23392 3290
rect 23444 3238 23456 3290
rect 23508 3238 23520 3290
rect 23572 3238 25852 3290
rect 1104 3216 25852 3238
rect 3050 3176 3056 3188
rect 1504 3148 3056 3176
rect 1504 3117 1532 3148
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 4580 3148 5733 3176
rect 4580 3136 4586 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 6822 3136 6828 3188
rect 6880 3136 6886 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 7156 3148 7205 3176
rect 7156 3136 7162 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 7282 3136 7288 3188
rect 7340 3136 7346 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 8938 3136 8944 3188
rect 8996 3176 9002 3188
rect 8996 3148 9996 3176
rect 8996 3136 9002 3148
rect 1489 3111 1547 3117
rect 1489 3077 1501 3111
rect 1535 3077 1547 3111
rect 1489 3071 1547 3077
rect 2590 3068 2596 3120
rect 2648 3068 2654 3120
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2774 3040 2780 3052
rect 2455 3012 2780 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 6012 3040 6040 3136
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6012 3012 6193 3040
rect 5905 3003 5963 3009
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6840 3040 6868 3136
rect 7300 3108 7328 3136
rect 8312 3108 8340 3136
rect 9766 3108 9772 3120
rect 7300 3080 7880 3108
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6840 3012 7389 3040
rect 6733 3003 6791 3009
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 3068 2972 3096 3003
rect 716 2944 3096 2972
rect 716 2932 722 2944
rect 5810 2932 5816 2984
rect 5868 2932 5874 2984
rect 5920 2972 5948 3003
rect 5920 2944 6408 2972
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 3237 2907 3295 2913
rect 2004 2876 2728 2904
rect 2004 2864 2010 2876
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 2700 2845 2728 2876
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 5442 2904 5448 2916
rect 3283 2876 5448 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 5828 2904 5856 2932
rect 6380 2913 6408 2944
rect 5997 2907 6055 2913
rect 5997 2904 6009 2907
rect 5828 2876 6009 2904
rect 5997 2873 6009 2876
rect 6043 2873 6055 2907
rect 5997 2867 6055 2873
rect 6365 2907 6423 2913
rect 6365 2873 6377 2907
rect 6411 2873 6423 2907
rect 6365 2867 6423 2873
rect 6546 2864 6552 2916
rect 6604 2904 6610 2916
rect 6748 2904 6776 3003
rect 7742 3000 7748 3052
rect 7800 3000 7806 3052
rect 6822 2932 6828 2984
rect 6880 2932 6886 2984
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7760 2972 7788 3000
rect 7055 2944 7788 2972
rect 7852 2972 7880 3080
rect 8036 3080 8340 3108
rect 9522 3080 9772 3108
rect 8036 3049 8064 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 9968 3108 9996 3148
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10778 3176 10784 3188
rect 10100 3148 10784 3176
rect 10100 3136 10106 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 12216 3148 13216 3176
rect 12216 3136 12222 3148
rect 10502 3108 10508 3120
rect 9968 3080 10508 3108
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 11790 3068 11796 3120
rect 11848 3068 11854 3120
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9640 3012 9873 3040
rect 9640 3000 9646 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 10137 3043 10195 3049
rect 10137 3040 10149 3043
rect 9861 3003 9919 3009
rect 10060 3012 10149 3040
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7852 2944 8309 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9766 2972 9772 2984
rect 9364 2944 9772 2972
rect 9364 2932 9370 2944
rect 9766 2932 9772 2944
rect 9824 2972 9830 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9824 2944 9965 2972
rect 9824 2932 9830 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 10060 2904 10088 3012
rect 10137 3009 10149 3012
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11296 3012 11529 3040
rect 11296 3000 11302 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 6604 2876 6868 2904
rect 6604 2864 6610 2876
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 72 2808 1593 2836
rect 72 2796 78 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2805 2743 2839
rect 6840 2836 6868 2876
rect 9324 2876 10088 2904
rect 10321 2907 10379 2913
rect 9324 2836 9352 2876
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 11514 2904 11520 2916
rect 10367 2876 11520 2904
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 12912 2904 12940 3026
rect 13188 2972 13216 3148
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 15562 3176 15568 3188
rect 14332 3148 15568 3176
rect 14332 3136 14338 3148
rect 15562 3136 15568 3148
rect 15620 3176 15626 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15620 3148 15669 3176
rect 15620 3136 15626 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 17221 3179 17279 3185
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 17402 3176 17408 3188
rect 17267 3148 17408 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 20898 3136 20904 3188
rect 20956 3136 20962 3188
rect 21821 3179 21879 3185
rect 21821 3145 21833 3179
rect 21867 3176 21879 3179
rect 22002 3176 22008 3188
rect 21867 3148 22008 3176
rect 21867 3145 21879 3148
rect 21821 3139 21879 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22189 3179 22247 3185
rect 22189 3145 22201 3179
rect 22235 3176 22247 3179
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 22235 3148 24409 3176
rect 22235 3145 22247 3148
rect 22189 3139 22247 3145
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 13280 3040 13308 3136
rect 14090 3068 14096 3120
rect 14148 3108 14154 3120
rect 14185 3111 14243 3117
rect 14185 3108 14197 3111
rect 14148 3080 14197 3108
rect 14148 3068 14154 3080
rect 14185 3077 14197 3080
rect 14231 3077 14243 3111
rect 14185 3071 14243 3077
rect 14918 3068 14924 3120
rect 14976 3068 14982 3120
rect 16669 3111 16727 3117
rect 16669 3077 16681 3111
rect 16715 3108 16727 3111
rect 17678 3108 17684 3120
rect 16715 3080 17684 3108
rect 16715 3077 16727 3080
rect 16669 3071 16727 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 21361 3111 21419 3117
rect 21361 3077 21373 3111
rect 21407 3108 21419 3111
rect 22094 3108 22100 3120
rect 21407 3080 22100 3108
rect 21407 3077 21419 3080
rect 21361 3071 21419 3077
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 22281 3111 22339 3117
rect 22281 3077 22293 3111
rect 22327 3108 22339 3111
rect 22830 3108 22836 3120
rect 22327 3080 22836 3108
rect 22327 3077 22339 3080
rect 22281 3071 22339 3077
rect 22830 3068 22836 3080
rect 22888 3068 22894 3120
rect 23106 3068 23112 3120
rect 23164 3108 23170 3120
rect 23164 3080 25268 3108
rect 23164 3068 23170 3080
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 13280 3012 13553 3040
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13906 3000 13912 3052
rect 13964 3000 13970 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17144 3012 17417 3040
rect 15470 2972 15476 2984
rect 13188 2944 15476 2972
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 17144 2981 17172 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 21266 3000 21272 3052
rect 21324 3000 21330 3052
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 21784 3012 22094 3040
rect 21784 3000 21790 3012
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 21048 2944 21465 2972
rect 21048 2932 21054 2944
rect 21453 2941 21465 2944
rect 21499 2941 21511 2975
rect 21453 2935 21511 2941
rect 13357 2907 13415 2913
rect 13357 2904 13369 2907
rect 12912 2876 13369 2904
rect 13357 2873 13369 2876
rect 13403 2873 13415 2907
rect 13357 2867 13415 2873
rect 17034 2864 17040 2916
rect 17092 2904 17098 2916
rect 17494 2904 17500 2916
rect 17092 2876 17500 2904
rect 17092 2864 17098 2876
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 22066 2904 22094 3012
rect 24578 3000 24584 3052
rect 24636 3000 24642 3052
rect 24670 3000 24676 3052
rect 24728 3040 24734 3052
rect 25240 3049 25268 3080
rect 24765 3043 24823 3049
rect 24765 3040 24777 3043
rect 24728 3012 24777 3040
rect 24728 3000 24734 3012
rect 24765 3009 24777 3012
rect 24811 3009 24823 3043
rect 24765 3003 24823 3009
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3009 25283 3043
rect 25225 3003 25283 3009
rect 22373 2975 22431 2981
rect 22373 2941 22385 2975
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 22388 2904 22416 2935
rect 22066 2876 22416 2904
rect 24670 2864 24676 2916
rect 24728 2904 24734 2916
rect 24728 2876 25452 2904
rect 24728 2864 24734 2876
rect 6840 2808 9352 2836
rect 2685 2799 2743 2805
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 9456 2808 9781 2836
rect 9456 2796 9462 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 10137 2839 10195 2845
rect 10137 2805 10149 2839
rect 10183 2836 10195 2839
rect 11330 2836 11336 2848
rect 10183 2808 11336 2836
rect 10183 2805 10195 2808
rect 10137 2799 10195 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 13262 2796 13268 2848
rect 13320 2796 13326 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 16850 2836 16856 2848
rect 15436 2808 16856 2836
rect 15436 2796 15442 2808
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 25041 2839 25099 2845
rect 25041 2805 25053 2839
rect 25087 2836 25099 2839
rect 25130 2836 25136 2848
rect 25087 2808 25136 2836
rect 25087 2805 25099 2808
rect 25041 2799 25099 2805
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 25424 2845 25452 2876
rect 25409 2839 25467 2845
rect 25409 2805 25421 2839
rect 25455 2805 25467 2839
rect 25409 2799 25467 2805
rect 1104 2746 25852 2768
rect 1104 2694 4043 2746
rect 4095 2694 4107 2746
rect 4159 2694 4171 2746
rect 4223 2694 4235 2746
rect 4287 2694 4299 2746
rect 4351 2694 10230 2746
rect 10282 2694 10294 2746
rect 10346 2694 10358 2746
rect 10410 2694 10422 2746
rect 10474 2694 10486 2746
rect 10538 2694 16417 2746
rect 16469 2694 16481 2746
rect 16533 2694 16545 2746
rect 16597 2694 16609 2746
rect 16661 2694 16673 2746
rect 16725 2694 22604 2746
rect 22656 2694 22668 2746
rect 22720 2694 22732 2746
rect 22784 2694 22796 2746
rect 22848 2694 22860 2746
rect 22912 2694 25852 2746
rect 1104 2672 25852 2694
rect 1302 2592 1308 2644
rect 1360 2632 1366 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 1360 2604 3157 2632
rect 1360 2592 1366 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 3145 2595 3203 2601
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 5166 2632 5172 2644
rect 4571 2604 5172 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 6546 2592 6552 2644
rect 6604 2592 6610 2644
rect 9122 2592 9128 2644
rect 9180 2592 9186 2644
rect 10594 2592 10600 2644
rect 10652 2592 10658 2644
rect 10778 2592 10784 2644
rect 10836 2592 10842 2644
rect 12526 2592 12532 2644
rect 12584 2592 12590 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 12860 2604 13645 2632
rect 12860 2592 12866 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 13814 2592 13820 2644
rect 13872 2592 13878 2644
rect 15013 2635 15071 2641
rect 15013 2601 15025 2635
rect 15059 2632 15071 2635
rect 15102 2632 15108 2644
rect 15059 2604 15108 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 17034 2592 17040 2644
rect 17092 2592 17098 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 21266 2632 21272 2644
rect 17267 2604 21272 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 21545 2635 21603 2641
rect 21545 2601 21557 2635
rect 21591 2632 21603 2635
rect 21910 2632 21916 2644
rect 21591 2604 21916 2632
rect 21591 2601 21603 2604
rect 21545 2595 21603 2601
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 8021 2567 8079 2573
rect 2516 2536 6914 2564
rect 2516 2437 2544 2536
rect 5442 2496 5448 2508
rect 3068 2468 5448 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2179 2400 2513 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 3068 2369 3096 2468
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 6886 2496 6914 2536
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 10796 2564 10824 2592
rect 13832 2564 13860 2592
rect 8067 2536 10824 2564
rect 12728 2536 13860 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 12434 2496 12440 2508
rect 6886 2468 12440 2496
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4120 2400 4353 2428
rect 4120 2388 4126 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9088 2400 9321 2428
rect 9088 2388 9094 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10134 2428 10140 2440
rect 9907 2400 10140 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 11054 2388 11060 2440
rect 11112 2388 11118 2440
rect 12250 2388 12256 2440
rect 12308 2388 12314 2440
rect 12728 2437 12756 2536
rect 13906 2524 13912 2576
rect 13964 2564 13970 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 13964 2536 14841 2564
rect 13964 2524 13970 2536
rect 14829 2533 14841 2536
rect 14875 2564 14887 2567
rect 17052 2564 17080 2592
rect 17770 2564 17776 2576
rect 14875 2536 17080 2564
rect 17604 2536 17776 2564
rect 14875 2533 14887 2536
rect 14829 2527 14887 2533
rect 15930 2496 15936 2508
rect 13096 2468 15936 2496
rect 13096 2437 13124 2468
rect 15930 2456 15936 2468
rect 15988 2496 15994 2508
rect 17604 2496 17632 2536
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 18966 2524 18972 2576
rect 19024 2564 19030 2576
rect 20257 2567 20315 2573
rect 20257 2564 20269 2567
rect 19024 2536 20269 2564
rect 19024 2524 19030 2536
rect 20257 2533 20269 2536
rect 20303 2533 20315 2567
rect 20257 2527 20315 2533
rect 20346 2524 20352 2576
rect 20404 2564 20410 2576
rect 24121 2567 24179 2573
rect 24121 2564 24133 2567
rect 20404 2536 24133 2564
rect 20404 2524 20410 2536
rect 24121 2533 24133 2536
rect 24167 2533 24179 2567
rect 24121 2527 24179 2533
rect 15988 2468 17632 2496
rect 15988 2456 15994 2468
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17736 2468 20392 2496
rect 17736 2456 17742 2468
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14550 2388 14556 2440
rect 14608 2388 14614 2440
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 15378 2388 15384 2440
rect 15436 2388 15442 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15528 2400 15884 2428
rect 15528 2388 15534 2400
rect 3053 2363 3111 2369
rect 1360 2332 2176 2360
rect 1360 2320 1366 2332
rect 2148 2292 2176 2332
rect 3053 2329 3065 2363
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 3878 2320 3884 2372
rect 3936 2320 3942 2372
rect 4709 2363 4767 2369
rect 4709 2329 4721 2363
rect 4755 2360 4767 2363
rect 5166 2360 5172 2372
rect 4755 2332 5172 2360
rect 4755 2329 4767 2332
rect 4709 2323 4767 2329
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 5350 2320 5356 2372
rect 5408 2320 5414 2372
rect 15396 2360 15424 2388
rect 11256 2332 15424 2360
rect 2593 2295 2651 2301
rect 2593 2292 2605 2295
rect 2148 2264 2605 2292
rect 2593 2261 2605 2264
rect 2639 2261 2651 2295
rect 2593 2255 2651 2261
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3476 2264 4169 2292
rect 3476 2252 3482 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4672 2264 4813 2292
rect 4672 2252 4678 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5629 2295 5687 2301
rect 5629 2292 5641 2295
rect 5316 2264 5641 2292
rect 5316 2252 5322 2264
rect 5629 2261 5641 2264
rect 5675 2261 5687 2295
rect 5629 2255 5687 2261
rect 7374 2252 7380 2304
rect 7432 2252 7438 2304
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 11256 2301 11284 2332
rect 15654 2320 15660 2372
rect 15712 2360 15718 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15712 2332 15761 2360
rect 15712 2320 15718 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15856 2360 15884 2400
rect 16758 2388 16764 2440
rect 16816 2388 16822 2440
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 16908 2400 17417 2428
rect 16908 2388 16914 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19576 2400 19809 2428
rect 19576 2388 19582 2400
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 18233 2363 18291 2369
rect 18233 2360 18245 2363
rect 15856 2332 18245 2360
rect 15749 2323 15807 2329
rect 18233 2329 18245 2332
rect 18279 2329 18291 2363
rect 18233 2323 18291 2329
rect 19334 2320 19340 2372
rect 19392 2320 19398 2372
rect 20364 2360 20392 2468
rect 20456 2468 21956 2496
rect 20456 2440 20484 2468
rect 20438 2388 20444 2440
rect 20496 2388 20502 2440
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 21726 2428 21732 2440
rect 21315 2400 21732 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 21726 2388 21732 2400
rect 21784 2388 21790 2440
rect 21928 2437 21956 2468
rect 21913 2431 21971 2437
rect 21913 2397 21925 2431
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 22922 2388 22928 2440
rect 22980 2388 22986 2440
rect 23934 2388 23940 2440
rect 23992 2388 23998 2440
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24912 2400 25145 2428
rect 24912 2388 24918 2400
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 24581 2363 24639 2369
rect 24581 2360 24593 2363
rect 20364 2332 24593 2360
rect 24581 2329 24593 2332
rect 24627 2329 24639 2363
rect 24581 2323 24639 2329
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 11241 2295 11299 2301
rect 11241 2261 11253 2295
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 12434 2252 12440 2304
rect 12492 2252 12498 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14976 2264 15301 2292
rect 14976 2252 14982 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15841 2295 15899 2301
rect 15841 2292 15853 2295
rect 15528 2264 15853 2292
rect 15528 2252 15534 2264
rect 15841 2261 15853 2264
rect 15887 2261 15899 2295
rect 15841 2255 15899 2261
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16540 2264 16865 2292
rect 16540 2252 16546 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18840 2264 19441 2292
rect 18840 2252 18846 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19978 2252 19984 2304
rect 20036 2252 20042 2304
rect 21726 2252 21732 2304
rect 21784 2292 21790 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21784 2264 22201 2292
rect 21784 2252 21790 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 24854 2252 24860 2304
rect 24912 2252 24918 2304
rect 25222 2252 25228 2304
rect 25280 2252 25286 2304
rect 1104 2202 25852 2224
rect 1104 2150 4703 2202
rect 4755 2150 4767 2202
rect 4819 2150 4831 2202
rect 4883 2150 4895 2202
rect 4947 2150 4959 2202
rect 5011 2150 10890 2202
rect 10942 2150 10954 2202
rect 11006 2150 11018 2202
rect 11070 2150 11082 2202
rect 11134 2150 11146 2202
rect 11198 2150 17077 2202
rect 17129 2150 17141 2202
rect 17193 2150 17205 2202
rect 17257 2150 17269 2202
rect 17321 2150 17333 2202
rect 17385 2150 23264 2202
rect 23316 2150 23328 2202
rect 23380 2150 23392 2202
rect 23444 2150 23456 2202
rect 23508 2150 23520 2202
rect 23572 2150 25852 2202
rect 1104 2128 25852 2150
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 5224 2060 6914 2088
rect 5224 2048 5230 2060
rect 5350 1980 5356 2032
rect 5408 1980 5414 2032
rect 5442 1980 5448 2032
rect 5500 1980 5506 2032
rect 6886 2020 6914 2060
rect 7374 2048 7380 2100
rect 7432 2088 7438 2100
rect 7432 2060 16574 2088
rect 7432 2048 7438 2060
rect 12710 2020 12716 2032
rect 6886 1992 12716 2020
rect 12710 1980 12716 1992
rect 12768 1980 12774 2032
rect 16546 2020 16574 2060
rect 22922 2048 22928 2100
rect 22980 2048 22986 2100
rect 22370 2020 22376 2032
rect 12820 1992 13032 2020
rect 16546 1992 22376 2020
rect 5368 1680 5396 1980
rect 5460 1748 5488 1980
rect 8110 1912 8116 1964
rect 8168 1952 8174 1964
rect 12820 1952 12848 1992
rect 8168 1924 12848 1952
rect 13004 1952 13032 1992
rect 22370 1980 22376 1992
rect 22428 1980 22434 2032
rect 19978 1952 19984 1964
rect 13004 1924 19984 1952
rect 8168 1912 8174 1924
rect 19978 1912 19984 1924
rect 20036 1912 20042 1964
rect 12618 1884 12624 1896
rect 9646 1856 12624 1884
rect 9646 1748 9674 1856
rect 12618 1844 12624 1856
rect 12676 1844 12682 1896
rect 12986 1844 12992 1896
rect 13044 1884 13050 1896
rect 19334 1884 19340 1896
rect 13044 1856 19340 1884
rect 13044 1844 13050 1856
rect 19334 1844 19340 1856
rect 19392 1844 19398 1896
rect 13446 1776 13452 1828
rect 13504 1816 13510 1828
rect 22940 1816 22968 2048
rect 13504 1788 22968 1816
rect 13504 1776 13510 1788
rect 5460 1720 9674 1748
rect 5368 1652 6914 1680
rect 6886 1544 6914 1652
rect 12434 1640 12440 1692
rect 12492 1680 12498 1692
rect 22462 1680 22468 1692
rect 12492 1652 22468 1680
rect 12492 1640 12498 1652
rect 22462 1640 22468 1652
rect 22520 1640 22526 1692
rect 13262 1544 13268 1556
rect 6886 1516 13268 1544
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 24578 1504 24584 1556
rect 24636 1544 24642 1556
rect 25774 1544 25780 1556
rect 24636 1516 25780 1544
rect 24636 1504 24642 1516
rect 25774 1504 25780 1516
rect 25832 1504 25838 1556
<< via1 >>
rect 4043 26630 4095 26682
rect 4107 26630 4159 26682
rect 4171 26630 4223 26682
rect 4235 26630 4287 26682
rect 4299 26630 4351 26682
rect 10230 26630 10282 26682
rect 10294 26630 10346 26682
rect 10358 26630 10410 26682
rect 10422 26630 10474 26682
rect 10486 26630 10538 26682
rect 16417 26630 16469 26682
rect 16481 26630 16533 26682
rect 16545 26630 16597 26682
rect 16609 26630 16661 26682
rect 16673 26630 16725 26682
rect 22604 26630 22656 26682
rect 22668 26630 22720 26682
rect 22732 26630 22784 26682
rect 22796 26630 22848 26682
rect 22860 26630 22912 26682
rect 1584 26571 1636 26580
rect 1584 26537 1593 26571
rect 1593 26537 1627 26571
rect 1627 26537 1636 26571
rect 1584 26528 1636 26537
rect 2228 26571 2280 26580
rect 2228 26537 2237 26571
rect 2237 26537 2271 26571
rect 2271 26537 2280 26571
rect 2228 26528 2280 26537
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 8392 26528 8444 26580
rect 11060 26571 11112 26580
rect 11060 26537 11069 26571
rect 11069 26537 11103 26571
rect 11103 26537 11112 26571
rect 11060 26528 11112 26537
rect 11612 26528 11664 26580
rect 14464 26571 14516 26580
rect 14464 26537 14473 26571
rect 14473 26537 14507 26571
rect 14507 26537 14516 26571
rect 14464 26528 14516 26537
rect 16764 26528 16816 26580
rect 5908 26460 5960 26512
rect 10692 26460 10744 26512
rect 17684 26528 17736 26580
rect 19064 26528 19116 26580
rect 19984 26528 20036 26580
rect 20720 26528 20772 26580
rect 23204 26528 23256 26580
rect 23940 26571 23992 26580
rect 23940 26537 23949 26571
rect 23949 26537 23983 26571
rect 23983 26537 23992 26571
rect 23940 26528 23992 26537
rect 18236 26460 18288 26512
rect 2688 26435 2740 26444
rect 2688 26401 2697 26435
rect 2697 26401 2731 26435
rect 2731 26401 2740 26435
rect 2688 26392 2740 26401
rect 1768 26256 1820 26308
rect 3240 26324 3292 26376
rect 5172 26324 5224 26376
rect 5816 26324 5868 26376
rect 6460 26324 6512 26376
rect 17960 26392 18012 26444
rect 22836 26460 22888 26512
rect 9312 26324 9364 26376
rect 9680 26324 9732 26376
rect 12256 26324 12308 26376
rect 12900 26324 12952 26376
rect 15476 26324 15528 26376
rect 3424 26256 3476 26308
rect 6828 26256 6880 26308
rect 7288 26299 7340 26308
rect 7288 26265 7297 26299
rect 7297 26265 7331 26299
rect 7331 26265 7340 26299
rect 7288 26256 7340 26265
rect 8208 26256 8260 26308
rect 10232 26256 10284 26308
rect 12072 26256 12124 26308
rect 14096 26256 14148 26308
rect 15016 26299 15068 26308
rect 15016 26265 15025 26299
rect 15025 26265 15059 26299
rect 15059 26265 15068 26299
rect 15016 26256 15068 26265
rect 15200 26256 15252 26308
rect 17408 26324 17460 26376
rect 18052 26324 18104 26376
rect 22100 26324 22152 26376
rect 16856 26256 16908 26308
rect 19432 26256 19484 26308
rect 21732 26256 21784 26308
rect 21916 26299 21968 26308
rect 21916 26265 21925 26299
rect 21925 26265 21959 26299
rect 21959 26265 21968 26299
rect 21916 26256 21968 26265
rect 24860 26460 24912 26512
rect 24584 26435 24636 26444
rect 24584 26401 24593 26435
rect 24593 26401 24627 26435
rect 24627 26401 24636 26435
rect 24584 26392 24636 26401
rect 25872 26324 25924 26376
rect 23848 26299 23900 26308
rect 23848 26265 23857 26299
rect 23857 26265 23891 26299
rect 23891 26265 23900 26299
rect 23848 26256 23900 26265
rect 5448 26231 5500 26240
rect 5448 26197 5457 26231
rect 5457 26197 5491 26231
rect 5491 26197 5500 26231
rect 5448 26188 5500 26197
rect 6092 26231 6144 26240
rect 6092 26197 6101 26231
rect 6101 26197 6135 26231
rect 6135 26197 6144 26231
rect 6092 26188 6144 26197
rect 6736 26231 6788 26240
rect 6736 26197 6745 26231
rect 6745 26197 6779 26231
rect 6779 26197 6788 26231
rect 6736 26188 6788 26197
rect 9680 26231 9732 26240
rect 9680 26197 9689 26231
rect 9689 26197 9723 26231
rect 9723 26197 9732 26231
rect 9680 26188 9732 26197
rect 12624 26188 12676 26240
rect 13176 26231 13228 26240
rect 13176 26197 13185 26231
rect 13185 26197 13219 26231
rect 13219 26197 13228 26231
rect 13176 26188 13228 26197
rect 14832 26188 14884 26240
rect 21272 26188 21324 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 23112 26188 23164 26240
rect 4703 26086 4755 26138
rect 4767 26086 4819 26138
rect 4831 26086 4883 26138
rect 4895 26086 4947 26138
rect 4959 26086 5011 26138
rect 10890 26086 10942 26138
rect 10954 26086 11006 26138
rect 11018 26086 11070 26138
rect 11082 26086 11134 26138
rect 11146 26086 11198 26138
rect 17077 26086 17129 26138
rect 17141 26086 17193 26138
rect 17205 26086 17257 26138
rect 17269 26086 17321 26138
rect 17333 26086 17385 26138
rect 23264 26086 23316 26138
rect 23328 26086 23380 26138
rect 23392 26086 23444 26138
rect 23456 26086 23508 26138
rect 23520 26086 23572 26138
rect 1032 25984 1084 26036
rect 5908 25984 5960 26036
rect 664 25916 716 25968
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 8576 25916 8628 25968
rect 9036 25916 9088 25968
rect 10140 25916 10192 25968
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 11980 25891 12032 25900
rect 11980 25857 11989 25891
rect 11989 25857 12023 25891
rect 12023 25857 12032 25891
rect 11980 25848 12032 25857
rect 8116 25823 8168 25832
rect 8116 25789 8125 25823
rect 8125 25789 8159 25823
rect 8159 25789 8168 25823
rect 8116 25780 8168 25789
rect 8300 25823 8352 25832
rect 8300 25789 8309 25823
rect 8309 25789 8343 25823
rect 8343 25789 8352 25823
rect 8300 25780 8352 25789
rect 8668 25780 8720 25832
rect 10876 25823 10928 25832
rect 10876 25789 10885 25823
rect 10885 25789 10919 25823
rect 10919 25789 10928 25823
rect 10876 25780 10928 25789
rect 20 25644 72 25696
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 3332 25687 3384 25696
rect 3332 25653 3341 25687
rect 3341 25653 3375 25687
rect 3375 25653 3384 25687
rect 3332 25644 3384 25653
rect 8576 25644 8628 25696
rect 8944 25644 8996 25696
rect 10600 25644 10652 25696
rect 11428 25712 11480 25764
rect 16212 25984 16264 26036
rect 23020 25984 23072 26036
rect 18788 25916 18840 25968
rect 15936 25848 15988 25900
rect 16120 25780 16172 25832
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 20352 25848 20404 25900
rect 22928 25848 22980 25900
rect 25320 25848 25372 25900
rect 26424 25848 26476 25900
rect 19708 25780 19760 25832
rect 11520 25687 11572 25696
rect 11520 25653 11529 25687
rect 11529 25653 11563 25687
rect 11563 25653 11572 25687
rect 11520 25644 11572 25653
rect 11796 25687 11848 25696
rect 11796 25653 11805 25687
rect 11805 25653 11839 25687
rect 11839 25653 11848 25687
rect 11796 25644 11848 25653
rect 18512 25644 18564 25696
rect 21548 25712 21600 25764
rect 24952 25823 25004 25832
rect 24952 25789 24961 25823
rect 24961 25789 24995 25823
rect 24995 25789 25004 25823
rect 24952 25780 25004 25789
rect 21180 25644 21232 25696
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 23940 25687 23992 25696
rect 23940 25653 23949 25687
rect 23949 25653 23983 25687
rect 23983 25653 23992 25687
rect 23940 25644 23992 25653
rect 4043 25542 4095 25594
rect 4107 25542 4159 25594
rect 4171 25542 4223 25594
rect 4235 25542 4287 25594
rect 4299 25542 4351 25594
rect 10230 25542 10282 25594
rect 10294 25542 10346 25594
rect 10358 25542 10410 25594
rect 10422 25542 10474 25594
rect 10486 25542 10538 25594
rect 16417 25542 16469 25594
rect 16481 25542 16533 25594
rect 16545 25542 16597 25594
rect 16609 25542 16661 25594
rect 16673 25542 16725 25594
rect 22604 25542 22656 25594
rect 22668 25542 22720 25594
rect 22732 25542 22784 25594
rect 22796 25542 22848 25594
rect 22860 25542 22912 25594
rect 1400 25440 1452 25492
rect 8208 25483 8260 25492
rect 8208 25449 8217 25483
rect 8217 25449 8251 25483
rect 8251 25449 8260 25483
rect 8208 25440 8260 25449
rect 9036 25440 9088 25492
rect 10140 25440 10192 25492
rect 8116 25372 8168 25424
rect 8300 25304 8352 25356
rect 11428 25440 11480 25492
rect 12900 25440 12952 25492
rect 12808 25372 12860 25424
rect 13820 25372 13872 25424
rect 15844 25483 15896 25492
rect 15844 25449 15853 25483
rect 15853 25449 15887 25483
rect 15887 25449 15896 25483
rect 15844 25440 15896 25449
rect 16856 25483 16908 25492
rect 16856 25449 16865 25483
rect 16865 25449 16899 25483
rect 16899 25449 16908 25483
rect 16856 25440 16908 25449
rect 17408 25483 17460 25492
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 17776 25440 17828 25492
rect 18788 25483 18840 25492
rect 18788 25449 18797 25483
rect 18797 25449 18831 25483
rect 18831 25449 18840 25483
rect 18788 25440 18840 25449
rect 19708 25440 19760 25492
rect 20352 25483 20404 25492
rect 20352 25449 20361 25483
rect 20361 25449 20395 25483
rect 20395 25449 20404 25483
rect 20352 25440 20404 25449
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 25504 25440 25556 25492
rect 20076 25372 20128 25424
rect 10416 25347 10468 25356
rect 1032 25236 1084 25288
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 2044 25168 2096 25220
rect 2688 25100 2740 25152
rect 8576 25236 8628 25288
rect 8944 25236 8996 25288
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 11520 25304 11572 25356
rect 13728 25304 13780 25356
rect 17868 25304 17920 25356
rect 18512 25347 18564 25356
rect 18512 25313 18521 25347
rect 18521 25313 18555 25347
rect 18555 25313 18564 25347
rect 18512 25304 18564 25313
rect 8576 25143 8628 25152
rect 8576 25109 8585 25143
rect 8585 25109 8619 25143
rect 8619 25109 8628 25143
rect 8576 25100 8628 25109
rect 9772 25168 9824 25220
rect 10508 25168 10560 25220
rect 10140 25143 10192 25152
rect 10140 25109 10149 25143
rect 10149 25109 10183 25143
rect 10183 25109 10192 25143
rect 10140 25100 10192 25109
rect 13176 25236 13228 25288
rect 11796 25168 11848 25220
rect 12716 25211 12768 25220
rect 12716 25177 12725 25211
rect 12725 25177 12759 25211
rect 12759 25177 12768 25211
rect 12716 25168 12768 25177
rect 14372 25211 14424 25220
rect 14372 25177 14381 25211
rect 14381 25177 14415 25211
rect 14415 25177 14424 25211
rect 14372 25168 14424 25177
rect 16672 25236 16724 25288
rect 11244 25100 11296 25152
rect 15108 25100 15160 25152
rect 16580 25100 16632 25152
rect 16856 25100 16908 25152
rect 16948 25100 17000 25152
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 19340 25236 19392 25288
rect 25780 25304 25832 25356
rect 24492 25236 24544 25288
rect 19524 25168 19576 25220
rect 17776 25143 17828 25152
rect 17776 25109 17785 25143
rect 17785 25109 17819 25143
rect 17819 25109 17828 25143
rect 17776 25100 17828 25109
rect 20996 25168 21048 25220
rect 21456 25168 21508 25220
rect 26148 25168 26200 25220
rect 22192 25143 22244 25152
rect 22192 25109 22201 25143
rect 22201 25109 22235 25143
rect 22235 25109 22244 25143
rect 22192 25100 22244 25109
rect 23756 25100 23808 25152
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 4703 24998 4755 25050
rect 4767 24998 4819 25050
rect 4831 24998 4883 25050
rect 4895 24998 4947 25050
rect 4959 24998 5011 25050
rect 10890 24998 10942 25050
rect 10954 24998 11006 25050
rect 11018 24998 11070 25050
rect 11082 24998 11134 25050
rect 11146 24998 11198 25050
rect 17077 24998 17129 25050
rect 17141 24998 17193 25050
rect 17205 24998 17257 25050
rect 17269 24998 17321 25050
rect 17333 24998 17385 25050
rect 23264 24998 23316 25050
rect 23328 24998 23380 25050
rect 23392 24998 23444 25050
rect 23456 24998 23508 25050
rect 23520 24998 23572 25050
rect 6368 24939 6420 24948
rect 6368 24905 6377 24939
rect 6377 24905 6411 24939
rect 6411 24905 6420 24939
rect 6368 24896 6420 24905
rect 11980 24939 12032 24948
rect 11980 24905 11989 24939
rect 11989 24905 12023 24939
rect 12023 24905 12032 24939
rect 11980 24896 12032 24905
rect 13176 24939 13228 24948
rect 13176 24905 13185 24939
rect 13185 24905 13219 24939
rect 13219 24905 13228 24939
rect 13176 24896 13228 24905
rect 14372 24896 14424 24948
rect 15292 24896 15344 24948
rect 16580 24896 16632 24948
rect 17408 24896 17460 24948
rect 19432 24896 19484 24948
rect 20996 24896 21048 24948
rect 6736 24871 6788 24880
rect 6736 24837 6745 24871
rect 6745 24837 6779 24871
rect 6779 24837 6788 24871
rect 6736 24828 6788 24837
rect 7656 24871 7708 24880
rect 7656 24837 7665 24871
rect 7665 24837 7699 24871
rect 7699 24837 7708 24871
rect 7656 24828 7708 24837
rect 8576 24828 8628 24880
rect 10784 24828 10836 24880
rect 12716 24871 12768 24880
rect 6828 24803 6880 24812
rect 6828 24769 6837 24803
rect 6837 24769 6871 24803
rect 6871 24769 6880 24803
rect 6828 24760 6880 24769
rect 8208 24803 8260 24812
rect 8208 24769 8217 24803
rect 8217 24769 8251 24803
rect 8251 24769 8260 24803
rect 8208 24760 8260 24769
rect 8300 24760 8352 24812
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 10600 24760 10652 24812
rect 12716 24837 12725 24871
rect 12725 24837 12759 24871
rect 12759 24837 12768 24871
rect 12716 24828 12768 24837
rect 14004 24828 14056 24880
rect 8116 24692 8168 24744
rect 10876 24735 10928 24744
rect 10876 24701 10885 24735
rect 10885 24701 10919 24735
rect 10919 24701 10928 24735
rect 10876 24692 10928 24701
rect 11980 24760 12032 24812
rect 12440 24803 12492 24812
rect 12440 24769 12449 24803
rect 12449 24769 12483 24803
rect 12483 24769 12492 24803
rect 12440 24760 12492 24769
rect 12164 24624 12216 24676
rect 12808 24624 12860 24676
rect 7288 24599 7340 24608
rect 7288 24565 7297 24599
rect 7297 24565 7331 24599
rect 7331 24565 7340 24599
rect 7288 24556 7340 24565
rect 9680 24556 9732 24608
rect 11336 24556 11388 24608
rect 11520 24556 11572 24608
rect 12256 24599 12308 24608
rect 12256 24565 12265 24599
rect 12265 24565 12299 24599
rect 12299 24565 12308 24599
rect 12256 24556 12308 24565
rect 13544 24735 13596 24744
rect 13544 24701 13553 24735
rect 13553 24701 13587 24735
rect 13587 24701 13596 24735
rect 13544 24692 13596 24701
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 16856 24828 16908 24880
rect 17592 24828 17644 24880
rect 17776 24828 17828 24880
rect 15108 24624 15160 24676
rect 13728 24556 13780 24608
rect 14648 24556 14700 24608
rect 16764 24760 16816 24812
rect 18144 24760 18196 24812
rect 21180 24828 21232 24880
rect 16212 24692 16264 24744
rect 16672 24624 16724 24676
rect 17316 24692 17368 24744
rect 15844 24556 15896 24608
rect 18144 24667 18196 24676
rect 18144 24633 18153 24667
rect 18153 24633 18187 24667
rect 18187 24633 18196 24667
rect 18144 24624 18196 24633
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 19616 24735 19668 24744
rect 19616 24701 19625 24735
rect 19625 24701 19659 24735
rect 19659 24701 19668 24735
rect 19616 24692 19668 24701
rect 21364 24803 21416 24812
rect 21364 24769 21373 24803
rect 21373 24769 21407 24803
rect 21407 24769 21416 24803
rect 21364 24760 21416 24769
rect 21088 24735 21140 24744
rect 21088 24701 21097 24735
rect 21097 24701 21131 24735
rect 21131 24701 21140 24735
rect 21088 24692 21140 24701
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 19800 24556 19852 24608
rect 4043 24454 4095 24506
rect 4107 24454 4159 24506
rect 4171 24454 4223 24506
rect 4235 24454 4287 24506
rect 4299 24454 4351 24506
rect 10230 24454 10282 24506
rect 10294 24454 10346 24506
rect 10358 24454 10410 24506
rect 10422 24454 10474 24506
rect 10486 24454 10538 24506
rect 16417 24454 16469 24506
rect 16481 24454 16533 24506
rect 16545 24454 16597 24506
rect 16609 24454 16661 24506
rect 16673 24454 16725 24506
rect 22604 24454 22656 24506
rect 22668 24454 22720 24506
rect 22732 24454 22784 24506
rect 22796 24454 22848 24506
rect 22860 24454 22912 24506
rect 7288 24352 7340 24404
rect 8668 24352 8720 24404
rect 10600 24352 10652 24404
rect 11428 24352 11480 24404
rect 12164 24352 12216 24404
rect 13544 24352 13596 24404
rect 8392 24148 8444 24200
rect 9128 24148 9180 24200
rect 940 24080 992 24132
rect 9772 24080 9824 24132
rect 11244 24216 11296 24268
rect 15568 24352 15620 24404
rect 15844 24352 15896 24404
rect 15936 24395 15988 24404
rect 15936 24361 15945 24395
rect 15945 24361 15979 24395
rect 15979 24361 15988 24395
rect 15936 24352 15988 24361
rect 16856 24352 16908 24404
rect 21364 24352 21416 24404
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 11336 24080 11388 24132
rect 12256 24080 12308 24132
rect 14648 24148 14700 24200
rect 15292 24148 15344 24200
rect 17132 24284 17184 24336
rect 20076 24327 20128 24336
rect 20076 24293 20085 24327
rect 20085 24293 20119 24327
rect 20119 24293 20128 24327
rect 20076 24284 20128 24293
rect 15660 24191 15712 24200
rect 15660 24157 15669 24191
rect 15669 24157 15703 24191
rect 15703 24157 15712 24191
rect 15660 24148 15712 24157
rect 16120 24148 16172 24200
rect 16948 24216 17000 24268
rect 17132 24148 17184 24200
rect 11520 24012 11572 24064
rect 14372 24012 14424 24064
rect 14464 24012 14516 24064
rect 15476 24012 15528 24064
rect 17408 24191 17460 24200
rect 17408 24157 17417 24191
rect 17417 24157 17451 24191
rect 17451 24157 17460 24191
rect 17408 24148 17460 24157
rect 17500 24148 17552 24200
rect 19524 24148 19576 24200
rect 19984 24148 20036 24200
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 18236 24080 18288 24132
rect 16212 24055 16264 24064
rect 16212 24021 16221 24055
rect 16221 24021 16255 24055
rect 16255 24021 16264 24055
rect 16212 24012 16264 24021
rect 16948 24012 17000 24064
rect 22008 24080 22060 24132
rect 21456 24055 21508 24064
rect 21456 24021 21465 24055
rect 21465 24021 21499 24055
rect 21499 24021 21508 24055
rect 21456 24012 21508 24021
rect 25412 24055 25464 24064
rect 25412 24021 25421 24055
rect 25421 24021 25455 24055
rect 25455 24021 25464 24055
rect 25412 24012 25464 24021
rect 4703 23910 4755 23962
rect 4767 23910 4819 23962
rect 4831 23910 4883 23962
rect 4895 23910 4947 23962
rect 4959 23910 5011 23962
rect 10890 23910 10942 23962
rect 10954 23910 11006 23962
rect 11018 23910 11070 23962
rect 11082 23910 11134 23962
rect 11146 23910 11198 23962
rect 17077 23910 17129 23962
rect 17141 23910 17193 23962
rect 17205 23910 17257 23962
rect 17269 23910 17321 23962
rect 17333 23910 17385 23962
rect 23264 23910 23316 23962
rect 23328 23910 23380 23962
rect 23392 23910 23444 23962
rect 23456 23910 23508 23962
rect 23520 23910 23572 23962
rect 1584 23808 1636 23860
rect 9634 23808 9686 23860
rect 9772 23808 9824 23860
rect 12440 23808 12492 23860
rect 14004 23808 14056 23860
rect 15660 23808 15712 23860
rect 15936 23808 15988 23860
rect 16304 23808 16356 23860
rect 19616 23808 19668 23860
rect 21364 23808 21416 23860
rect 21456 23808 21508 23860
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 11796 23783 11848 23792
rect 11796 23749 11805 23783
rect 11805 23749 11839 23783
rect 11839 23749 11848 23783
rect 11796 23740 11848 23749
rect 11980 23740 12032 23792
rect 13820 23740 13872 23792
rect 5264 23672 5316 23724
rect 6184 23672 6236 23724
rect 5724 23604 5776 23656
rect 6000 23604 6052 23656
rect 1584 23579 1636 23588
rect 1584 23545 1593 23579
rect 1593 23545 1627 23579
rect 1627 23545 1636 23579
rect 1584 23536 1636 23545
rect 5908 23536 5960 23588
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 9496 23672 9548 23724
rect 9772 23715 9824 23724
rect 9772 23681 9781 23715
rect 9781 23681 9815 23715
rect 9815 23681 9824 23715
rect 9772 23672 9824 23681
rect 10140 23604 10192 23656
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 10508 23604 10560 23656
rect 15660 23672 15712 23724
rect 16028 23715 16080 23724
rect 16028 23681 16043 23715
rect 16043 23681 16077 23715
rect 16077 23681 16080 23715
rect 16028 23672 16080 23681
rect 10048 23536 10100 23588
rect 10416 23536 10468 23588
rect 12256 23536 12308 23588
rect 12808 23536 12860 23588
rect 16028 23536 16080 23588
rect 16764 23740 16816 23792
rect 19340 23740 19392 23792
rect 17592 23672 17644 23724
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 20720 23715 20772 23724
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 22008 23740 22060 23792
rect 20904 23604 20956 23656
rect 16396 23536 16448 23588
rect 19524 23536 19576 23588
rect 21548 23647 21600 23656
rect 21548 23613 21557 23647
rect 21557 23613 21591 23647
rect 21591 23613 21600 23647
rect 21548 23604 21600 23613
rect 22192 23604 22244 23656
rect 25596 23604 25648 23656
rect 5540 23468 5592 23520
rect 6828 23468 6880 23520
rect 8668 23468 8720 23520
rect 9772 23468 9824 23520
rect 9956 23468 10008 23520
rect 16948 23468 17000 23520
rect 20996 23468 21048 23520
rect 21548 23468 21600 23520
rect 21824 23468 21876 23520
rect 23756 23468 23808 23520
rect 24308 23468 24360 23520
rect 25504 23511 25556 23520
rect 25504 23477 25513 23511
rect 25513 23477 25547 23511
rect 25547 23477 25556 23511
rect 25504 23468 25556 23477
rect 25780 23468 25832 23520
rect 4043 23366 4095 23418
rect 4107 23366 4159 23418
rect 4171 23366 4223 23418
rect 4235 23366 4287 23418
rect 4299 23366 4351 23418
rect 10230 23366 10282 23418
rect 10294 23366 10346 23418
rect 10358 23366 10410 23418
rect 10422 23366 10474 23418
rect 10486 23366 10538 23418
rect 16417 23366 16469 23418
rect 16481 23366 16533 23418
rect 16545 23366 16597 23418
rect 16609 23366 16661 23418
rect 16673 23366 16725 23418
rect 22604 23366 22656 23418
rect 22668 23366 22720 23418
rect 22732 23366 22784 23418
rect 22796 23366 22848 23418
rect 22860 23366 22912 23418
rect 6828 23264 6880 23316
rect 3608 23196 3660 23248
rect 5540 23103 5592 23112
rect 5540 23069 5552 23103
rect 5552 23069 5586 23103
rect 5586 23069 5592 23103
rect 5540 23060 5592 23069
rect 5724 23060 5776 23112
rect 5816 23103 5868 23112
rect 5816 23069 5825 23103
rect 5825 23069 5859 23103
rect 5859 23069 5868 23103
rect 5816 23060 5868 23069
rect 5908 23103 5960 23112
rect 5908 23069 5917 23103
rect 5917 23069 5951 23103
rect 5951 23069 5960 23103
rect 5908 23060 5960 23069
rect 6368 23171 6420 23180
rect 6368 23137 6377 23171
rect 6377 23137 6411 23171
rect 6411 23137 6420 23171
rect 6368 23128 6420 23137
rect 6644 23171 6696 23180
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 7564 23128 7616 23180
rect 8852 23128 8904 23180
rect 9772 23264 9824 23316
rect 14464 23264 14516 23316
rect 15660 23264 15712 23316
rect 15936 23264 15988 23316
rect 16948 23264 17000 23316
rect 20720 23264 20772 23316
rect 20904 23307 20956 23316
rect 20904 23273 20913 23307
rect 20913 23273 20947 23307
rect 20947 23273 20956 23307
rect 20904 23264 20956 23273
rect 16212 23196 16264 23248
rect 9588 23128 9640 23180
rect 6092 23060 6144 23112
rect 7656 23060 7708 23112
rect 6184 22992 6236 23044
rect 9220 23035 9272 23044
rect 9220 23001 9229 23035
rect 9229 23001 9263 23035
rect 9263 23001 9272 23035
rect 9220 22992 9272 23001
rect 9956 22992 10008 23044
rect 11336 22992 11388 23044
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 14556 23060 14608 23112
rect 16120 23060 16172 23112
rect 16304 23060 16356 23112
rect 16764 23060 16816 23112
rect 19524 23239 19576 23248
rect 19524 23205 19533 23239
rect 19533 23205 19567 23239
rect 19567 23205 19576 23239
rect 19524 23196 19576 23205
rect 20076 23196 20128 23248
rect 19984 23128 20036 23180
rect 17408 23060 17460 23112
rect 4620 22924 4672 22976
rect 5264 22967 5316 22976
rect 5264 22933 5273 22967
rect 5273 22933 5307 22967
rect 5307 22933 5316 22967
rect 5264 22924 5316 22933
rect 6828 22924 6880 22976
rect 7104 22967 7156 22976
rect 7104 22933 7113 22967
rect 7113 22933 7147 22967
rect 7147 22933 7156 22967
rect 7104 22924 7156 22933
rect 7288 22967 7340 22976
rect 7288 22933 7297 22967
rect 7297 22933 7331 22967
rect 7331 22933 7340 22967
rect 7288 22924 7340 22933
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 16304 22924 16356 22976
rect 17500 22924 17552 22976
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 20628 23128 20680 23180
rect 21916 23128 21968 23180
rect 20536 23103 20588 23112
rect 20536 23069 20545 23103
rect 20545 23069 20579 23103
rect 20579 23069 20588 23103
rect 20536 23060 20588 23069
rect 21272 22967 21324 22976
rect 21272 22933 21281 22967
rect 21281 22933 21315 22967
rect 21315 22933 21324 22967
rect 21272 22924 21324 22933
rect 4703 22822 4755 22874
rect 4767 22822 4819 22874
rect 4831 22822 4883 22874
rect 4895 22822 4947 22874
rect 4959 22822 5011 22874
rect 10890 22822 10942 22874
rect 10954 22822 11006 22874
rect 11018 22822 11070 22874
rect 11082 22822 11134 22874
rect 11146 22822 11198 22874
rect 17077 22822 17129 22874
rect 17141 22822 17193 22874
rect 17205 22822 17257 22874
rect 17269 22822 17321 22874
rect 17333 22822 17385 22874
rect 23264 22822 23316 22874
rect 23328 22822 23380 22874
rect 23392 22822 23444 22874
rect 23456 22822 23508 22874
rect 23520 22822 23572 22874
rect 3056 22720 3108 22772
rect 3700 22720 3752 22772
rect 5724 22720 5776 22772
rect 6644 22720 6696 22772
rect 3792 22652 3844 22704
rect 2504 22584 2556 22636
rect 7012 22652 7064 22704
rect 8208 22720 8260 22772
rect 9220 22720 9272 22772
rect 10140 22720 10192 22772
rect 11336 22720 11388 22772
rect 12164 22720 12216 22772
rect 12624 22720 12676 22772
rect 14188 22763 14240 22772
rect 14188 22729 14197 22763
rect 14197 22729 14231 22763
rect 14231 22729 14240 22763
rect 14188 22720 14240 22729
rect 14280 22720 14332 22772
rect 5080 22627 5132 22636
rect 5080 22593 5089 22627
rect 5089 22593 5123 22627
rect 5123 22593 5132 22627
rect 5080 22584 5132 22593
rect 7196 22584 7248 22636
rect 3608 22516 3660 22568
rect 5540 22516 5592 22568
rect 5724 22516 5776 22568
rect 6184 22516 6236 22568
rect 6920 22516 6972 22568
rect 7564 22516 7616 22568
rect 12348 22652 12400 22704
rect 8024 22627 8076 22636
rect 8024 22593 8033 22627
rect 8033 22593 8067 22627
rect 8067 22593 8076 22627
rect 8024 22584 8076 22593
rect 4436 22448 4488 22500
rect 11244 22584 11296 22636
rect 9680 22516 9732 22568
rect 13636 22559 13688 22568
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 15660 22652 15712 22704
rect 940 22380 992 22432
rect 2228 22380 2280 22432
rect 4528 22423 4580 22432
rect 4528 22389 4537 22423
rect 4537 22389 4571 22423
rect 4571 22389 4580 22423
rect 4528 22380 4580 22389
rect 8208 22448 8260 22500
rect 8944 22380 8996 22432
rect 10140 22491 10192 22500
rect 10140 22457 10149 22491
rect 10149 22457 10183 22491
rect 10183 22457 10192 22491
rect 10140 22448 10192 22457
rect 14556 22516 14608 22568
rect 15936 22584 15988 22636
rect 15752 22516 15804 22568
rect 17316 22720 17368 22772
rect 17408 22720 17460 22772
rect 19708 22720 19760 22772
rect 21916 22720 21968 22772
rect 17500 22652 17552 22704
rect 16212 22559 16264 22568
rect 16212 22525 16221 22559
rect 16221 22525 16255 22559
rect 16255 22525 16264 22559
rect 16212 22516 16264 22525
rect 14188 22448 14240 22500
rect 13636 22380 13688 22432
rect 16212 22380 16264 22432
rect 17776 22584 17828 22636
rect 19340 22584 19392 22636
rect 20996 22652 21048 22704
rect 17316 22559 17368 22568
rect 17316 22525 17325 22559
rect 17325 22525 17359 22559
rect 17359 22525 17368 22559
rect 17316 22516 17368 22525
rect 17592 22516 17644 22568
rect 20720 22516 20772 22568
rect 25964 22516 26016 22568
rect 17408 22448 17460 22500
rect 16948 22380 17000 22432
rect 18052 22380 18104 22432
rect 19984 22380 20036 22432
rect 26240 22380 26292 22432
rect 4043 22278 4095 22330
rect 4107 22278 4159 22330
rect 4171 22278 4223 22330
rect 4235 22278 4287 22330
rect 4299 22278 4351 22330
rect 10230 22278 10282 22330
rect 10294 22278 10346 22330
rect 10358 22278 10410 22330
rect 10422 22278 10474 22330
rect 10486 22278 10538 22330
rect 16417 22278 16469 22330
rect 16481 22278 16533 22330
rect 16545 22278 16597 22330
rect 16609 22278 16661 22330
rect 16673 22278 16725 22330
rect 22604 22278 22656 22330
rect 22668 22278 22720 22330
rect 22732 22278 22784 22330
rect 22796 22278 22848 22330
rect 22860 22278 22912 22330
rect 2228 22176 2280 22228
rect 3608 22219 3660 22228
rect 3608 22185 3617 22219
rect 3617 22185 3651 22219
rect 3651 22185 3660 22219
rect 3608 22176 3660 22185
rect 3792 22219 3844 22228
rect 3792 22185 3801 22219
rect 3801 22185 3835 22219
rect 3835 22185 3844 22219
rect 3792 22176 3844 22185
rect 4436 22176 4488 22228
rect 5816 22176 5868 22228
rect 6920 22176 6972 22228
rect 7288 22176 7340 22228
rect 7564 22176 7616 22228
rect 10232 22176 10284 22228
rect 12256 22176 12308 22228
rect 12348 22219 12400 22228
rect 12348 22185 12357 22219
rect 12357 22185 12391 22219
rect 12391 22185 12400 22219
rect 12348 22176 12400 22185
rect 12900 22176 12952 22228
rect 13636 22176 13688 22228
rect 14096 22176 14148 22228
rect 15936 22219 15988 22228
rect 15936 22185 15945 22219
rect 15945 22185 15979 22219
rect 15979 22185 15988 22219
rect 15936 22176 15988 22185
rect 16304 22176 16356 22228
rect 5356 22108 5408 22160
rect 2136 21904 2188 21956
rect 4436 21904 4488 21956
rect 5172 21904 5224 21956
rect 5816 21972 5868 22024
rect 2412 21836 2464 21888
rect 5632 21836 5684 21888
rect 5724 21836 5776 21888
rect 5908 21879 5960 21888
rect 5908 21845 5917 21879
rect 5917 21845 5951 21879
rect 5951 21845 5960 21879
rect 5908 21836 5960 21845
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6644 21972 6696 21981
rect 6828 21972 6880 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 8300 21972 8352 22024
rect 8668 22108 8720 22160
rect 15660 22108 15712 22160
rect 10140 22040 10192 22092
rect 11612 22040 11664 22092
rect 12164 22040 12216 22092
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 8852 21972 8904 22024
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 10784 21972 10836 22024
rect 6552 21836 6604 21888
rect 9588 21836 9640 21888
rect 10784 21836 10836 21888
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11336 21972 11388 21981
rect 11796 22015 11848 22024
rect 11796 21981 11805 22015
rect 11805 21981 11839 22015
rect 11839 21981 11848 22015
rect 11796 21972 11848 21981
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 17316 22176 17368 22228
rect 17684 22176 17736 22228
rect 17868 22176 17920 22228
rect 13728 21972 13780 22024
rect 16212 21972 16264 22024
rect 16764 22015 16816 22024
rect 16764 21981 16773 22015
rect 16773 21981 16807 22015
rect 16807 21981 16816 22015
rect 16764 21972 16816 21981
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 17408 21972 17460 22024
rect 17592 21972 17644 22024
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 20720 22176 20772 22228
rect 20628 22108 20680 22160
rect 19248 22083 19300 22092
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 11428 21904 11480 21956
rect 13636 21904 13688 21956
rect 13084 21836 13136 21888
rect 13176 21879 13228 21888
rect 13176 21845 13185 21879
rect 13185 21845 13219 21879
rect 13219 21845 13228 21879
rect 13176 21836 13228 21845
rect 13820 21836 13872 21888
rect 14464 21836 14516 21888
rect 16856 21836 16908 21888
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 19524 21947 19576 21956
rect 19524 21913 19533 21947
rect 19533 21913 19567 21947
rect 19567 21913 19576 21947
rect 19524 21904 19576 21913
rect 19984 21904 20036 21956
rect 25964 21904 26016 21956
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 18972 21836 19024 21888
rect 20536 21836 20588 21888
rect 4703 21734 4755 21786
rect 4767 21734 4819 21786
rect 4831 21734 4883 21786
rect 4895 21734 4947 21786
rect 4959 21734 5011 21786
rect 10890 21734 10942 21786
rect 10954 21734 11006 21786
rect 11018 21734 11070 21786
rect 11082 21734 11134 21786
rect 11146 21734 11198 21786
rect 17077 21734 17129 21786
rect 17141 21734 17193 21786
rect 17205 21734 17257 21786
rect 17269 21734 17321 21786
rect 17333 21734 17385 21786
rect 23264 21734 23316 21786
rect 23328 21734 23380 21786
rect 23392 21734 23444 21786
rect 23456 21734 23508 21786
rect 23520 21734 23572 21786
rect 2136 21675 2188 21684
rect 2136 21641 2145 21675
rect 2145 21641 2179 21675
rect 2179 21641 2188 21675
rect 2136 21632 2188 21641
rect 2412 21632 2464 21684
rect 8392 21632 8444 21684
rect 8852 21632 8904 21684
rect 11336 21632 11388 21684
rect 13176 21632 13228 21684
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 3332 21564 3384 21616
rect 4528 21564 4580 21616
rect 5632 21564 5684 21616
rect 6000 21564 6052 21616
rect 6368 21607 6420 21616
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 5264 21496 5316 21548
rect 6092 21539 6144 21548
rect 6092 21505 6101 21539
rect 6101 21505 6135 21539
rect 6135 21505 6144 21539
rect 6092 21496 6144 21505
rect 6368 21573 6377 21607
rect 6377 21573 6411 21607
rect 6411 21573 6420 21607
rect 6368 21564 6420 21573
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 5172 21471 5224 21480
rect 5172 21437 5181 21471
rect 5181 21437 5215 21471
rect 5215 21437 5224 21471
rect 5172 21428 5224 21437
rect 5724 21428 5776 21480
rect 6644 21471 6696 21480
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 940 21292 992 21344
rect 5540 21403 5592 21412
rect 5540 21369 5549 21403
rect 5549 21369 5583 21403
rect 5583 21369 5592 21403
rect 5540 21360 5592 21369
rect 5816 21360 5868 21412
rect 7104 21607 7156 21616
rect 7104 21573 7113 21607
rect 7113 21573 7147 21607
rect 7147 21573 7156 21607
rect 7104 21564 7156 21573
rect 7196 21564 7248 21616
rect 7656 21564 7708 21616
rect 9956 21564 10008 21616
rect 10784 21564 10836 21616
rect 7104 21428 7156 21480
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 9588 21496 9640 21548
rect 12256 21496 12308 21548
rect 13728 21564 13780 21616
rect 16212 21632 16264 21684
rect 16764 21632 16816 21684
rect 16672 21607 16724 21616
rect 16672 21573 16681 21607
rect 16681 21573 16715 21607
rect 16715 21573 16724 21607
rect 19524 21632 19576 21684
rect 21272 21632 21324 21684
rect 16672 21564 16724 21573
rect 16948 21496 17000 21548
rect 17224 21496 17276 21548
rect 25228 21564 25280 21616
rect 18328 21496 18380 21548
rect 20168 21496 20220 21548
rect 21640 21539 21692 21548
rect 21640 21505 21649 21539
rect 21649 21505 21683 21539
rect 21683 21505 21692 21539
rect 21640 21496 21692 21505
rect 21824 21496 21876 21548
rect 9680 21428 9732 21480
rect 4988 21292 5040 21344
rect 7564 21360 7616 21412
rect 12808 21428 12860 21480
rect 14188 21428 14240 21480
rect 10140 21292 10192 21344
rect 15476 21360 15528 21412
rect 16948 21360 17000 21412
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 18052 21428 18104 21480
rect 19432 21428 19484 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 20628 21471 20680 21480
rect 20628 21437 20637 21471
rect 20637 21437 20671 21471
rect 20671 21437 20680 21471
rect 20628 21428 20680 21437
rect 17592 21360 17644 21412
rect 17684 21403 17736 21412
rect 17684 21369 17693 21403
rect 17693 21369 17727 21403
rect 17727 21369 17736 21403
rect 17684 21360 17736 21369
rect 20260 21360 20312 21412
rect 13084 21292 13136 21344
rect 24124 21471 24176 21480
rect 24124 21437 24133 21471
rect 24133 21437 24167 21471
rect 24167 21437 24176 21471
rect 24124 21428 24176 21437
rect 21456 21335 21508 21344
rect 21456 21301 21465 21335
rect 21465 21301 21499 21335
rect 21499 21301 21508 21335
rect 21456 21292 21508 21301
rect 23664 21292 23716 21344
rect 4043 21190 4095 21242
rect 4107 21190 4159 21242
rect 4171 21190 4223 21242
rect 4235 21190 4287 21242
rect 4299 21190 4351 21242
rect 10230 21190 10282 21242
rect 10294 21190 10346 21242
rect 10358 21190 10410 21242
rect 10422 21190 10474 21242
rect 10486 21190 10538 21242
rect 16417 21190 16469 21242
rect 16481 21190 16533 21242
rect 16545 21190 16597 21242
rect 16609 21190 16661 21242
rect 16673 21190 16725 21242
rect 22604 21190 22656 21242
rect 22668 21190 22720 21242
rect 22732 21190 22784 21242
rect 22796 21190 22848 21242
rect 22860 21190 22912 21242
rect 2320 21088 2372 21140
rect 3240 21088 3292 21140
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 5540 21088 5592 21140
rect 6552 21088 6604 21140
rect 7288 21088 7340 21140
rect 5908 21020 5960 21072
rect 7104 21020 7156 21072
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 4436 20952 4488 21004
rect 10140 21020 10192 21072
rect 11428 21088 11480 21140
rect 11612 21131 11664 21140
rect 11612 21097 11621 21131
rect 11621 21097 11655 21131
rect 11655 21097 11664 21131
rect 11612 21088 11664 21097
rect 11796 21020 11848 21072
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 13728 21088 13780 21140
rect 19340 21088 19392 21140
rect 21640 21088 21692 21140
rect 7840 20952 7892 21004
rect 20628 21063 20680 21072
rect 20628 21029 20637 21063
rect 20637 21029 20671 21063
rect 20671 21029 20680 21063
rect 20628 21020 20680 21029
rect 26332 21020 26384 21072
rect 5172 20927 5224 20936
rect 5172 20893 5181 20927
rect 5181 20893 5215 20927
rect 5215 20893 5224 20927
rect 5172 20884 5224 20893
rect 5264 20884 5316 20936
rect 5540 20884 5592 20936
rect 8300 20884 8352 20936
rect 2964 20816 3016 20868
rect 4988 20816 5040 20868
rect 7564 20816 7616 20868
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 10324 20884 10376 20936
rect 9680 20859 9732 20868
rect 9680 20825 9689 20859
rect 9689 20825 9723 20859
rect 9723 20825 9732 20859
rect 9680 20816 9732 20825
rect 11428 20884 11480 20936
rect 13820 20927 13872 20936
rect 13820 20893 13829 20927
rect 13829 20893 13863 20927
rect 13863 20893 13872 20927
rect 13820 20884 13872 20893
rect 14188 20884 14240 20936
rect 14372 20884 14424 20936
rect 14464 20927 14516 20936
rect 14464 20893 14473 20927
rect 14473 20893 14507 20927
rect 14507 20893 14516 20927
rect 14464 20884 14516 20893
rect 11244 20816 11296 20868
rect 11520 20859 11572 20868
rect 11520 20825 11529 20859
rect 11529 20825 11563 20859
rect 11563 20825 11572 20859
rect 11520 20816 11572 20825
rect 11888 20859 11940 20868
rect 11888 20825 11897 20859
rect 11897 20825 11931 20859
rect 11931 20825 11940 20859
rect 11888 20816 11940 20825
rect 13176 20816 13228 20868
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 6644 20748 6696 20800
rect 7380 20748 7432 20800
rect 8576 20791 8628 20800
rect 8576 20757 8585 20791
rect 8585 20757 8619 20791
rect 8619 20757 8628 20791
rect 8576 20748 8628 20757
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 10140 20791 10192 20800
rect 10140 20757 10149 20791
rect 10149 20757 10183 20791
rect 10183 20757 10192 20791
rect 10140 20748 10192 20757
rect 10324 20748 10376 20800
rect 12992 20748 13044 20800
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 14740 20884 14792 20936
rect 24952 20952 25004 21004
rect 16212 20884 16264 20936
rect 20536 20884 20588 20936
rect 14280 20748 14332 20800
rect 19340 20816 19392 20868
rect 21180 20859 21232 20868
rect 21180 20825 21189 20859
rect 21189 20825 21223 20859
rect 21223 20825 21232 20859
rect 21180 20816 21232 20825
rect 21456 20816 21508 20868
rect 17408 20748 17460 20800
rect 22192 20748 22244 20800
rect 4703 20646 4755 20698
rect 4767 20646 4819 20698
rect 4831 20646 4883 20698
rect 4895 20646 4947 20698
rect 4959 20646 5011 20698
rect 10890 20646 10942 20698
rect 10954 20646 11006 20698
rect 11018 20646 11070 20698
rect 11082 20646 11134 20698
rect 11146 20646 11198 20698
rect 17077 20646 17129 20698
rect 17141 20646 17193 20698
rect 17205 20646 17257 20698
rect 17269 20646 17321 20698
rect 17333 20646 17385 20698
rect 23264 20646 23316 20698
rect 23328 20646 23380 20698
rect 23392 20646 23444 20698
rect 23456 20646 23508 20698
rect 23520 20646 23572 20698
rect 25964 20680 26016 20732
rect 4804 20544 4856 20596
rect 3240 20476 3292 20528
rect 9588 20544 9640 20596
rect 10140 20544 10192 20596
rect 2964 20383 3016 20392
rect 2964 20349 2973 20383
rect 2973 20349 3007 20383
rect 3007 20349 3016 20383
rect 2964 20340 3016 20349
rect 3792 20408 3844 20460
rect 9956 20476 10008 20528
rect 7104 20340 7156 20392
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 11152 20408 11204 20460
rect 8668 20340 8720 20392
rect 9312 20340 9364 20392
rect 11888 20544 11940 20596
rect 12716 20544 12768 20596
rect 12808 20587 12860 20596
rect 12808 20553 12817 20587
rect 12817 20553 12851 20587
rect 12851 20553 12860 20587
rect 12808 20544 12860 20553
rect 13176 20544 13228 20596
rect 21180 20544 21232 20596
rect 11520 20451 11572 20460
rect 11520 20417 11529 20451
rect 11529 20417 11563 20451
rect 11563 20417 11572 20451
rect 11520 20408 11572 20417
rect 11888 20408 11940 20460
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 16120 20476 16172 20528
rect 3240 20315 3292 20324
rect 3240 20281 3249 20315
rect 3249 20281 3283 20315
rect 3283 20281 3292 20315
rect 3240 20272 3292 20281
rect 3516 20247 3568 20256
rect 3516 20213 3525 20247
rect 3525 20213 3559 20247
rect 3559 20213 3568 20247
rect 3516 20204 3568 20213
rect 3608 20204 3660 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 8392 20204 8444 20256
rect 8852 20204 8904 20256
rect 12532 20340 12584 20392
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 15936 20408 15988 20460
rect 16304 20408 16356 20460
rect 18328 20340 18380 20392
rect 20444 20408 20496 20460
rect 22192 20544 22244 20596
rect 23664 20544 23716 20596
rect 22468 20408 22520 20460
rect 23112 20408 23164 20460
rect 19800 20340 19852 20392
rect 9956 20272 10008 20324
rect 11428 20272 11480 20324
rect 12256 20272 12308 20324
rect 15384 20272 15436 20324
rect 15936 20272 15988 20324
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 11336 20204 11388 20256
rect 11704 20247 11756 20256
rect 11704 20213 11713 20247
rect 11713 20213 11747 20247
rect 11747 20213 11756 20247
rect 11704 20204 11756 20213
rect 12440 20204 12492 20256
rect 18604 20247 18656 20256
rect 18604 20213 18613 20247
rect 18613 20213 18647 20247
rect 18647 20213 18656 20247
rect 18604 20204 18656 20213
rect 20076 20204 20128 20256
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 22192 20204 22244 20256
rect 23664 20204 23716 20256
rect 4043 20102 4095 20154
rect 4107 20102 4159 20154
rect 4171 20102 4223 20154
rect 4235 20102 4287 20154
rect 4299 20102 4351 20154
rect 10230 20102 10282 20154
rect 10294 20102 10346 20154
rect 10358 20102 10410 20154
rect 10422 20102 10474 20154
rect 10486 20102 10538 20154
rect 16417 20102 16469 20154
rect 16481 20102 16533 20154
rect 16545 20102 16597 20154
rect 16609 20102 16661 20154
rect 16673 20102 16725 20154
rect 22604 20102 22656 20154
rect 22668 20102 22720 20154
rect 22732 20102 22784 20154
rect 22796 20102 22848 20154
rect 22860 20102 22912 20154
rect 2596 20000 2648 20052
rect 4068 20000 4120 20052
rect 4712 20000 4764 20052
rect 6644 20000 6696 20052
rect 7288 20000 7340 20052
rect 7656 20000 7708 20052
rect 8392 20000 8444 20052
rect 9036 20000 9088 20052
rect 9220 20000 9272 20052
rect 9680 20000 9732 20052
rect 10140 20000 10192 20052
rect 11152 20000 11204 20052
rect 11520 20000 11572 20052
rect 12440 20000 12492 20052
rect 12532 20000 12584 20052
rect 14188 20000 14240 20052
rect 14648 20000 14700 20052
rect 15384 20000 15436 20052
rect 1676 19864 1728 19916
rect 2688 19864 2740 19916
rect 3700 19864 3752 19916
rect 4068 19864 4120 19916
rect 4252 19864 4304 19916
rect 4804 19864 4856 19916
rect 6828 19975 6880 19984
rect 6828 19941 6837 19975
rect 6837 19941 6871 19975
rect 6871 19941 6880 19975
rect 6828 19932 6880 19941
rect 7104 19932 7156 19984
rect 11336 19932 11388 19984
rect 4436 19796 4488 19848
rect 4528 19796 4580 19848
rect 2044 19771 2096 19780
rect 2044 19737 2053 19771
rect 2053 19737 2087 19771
rect 2087 19737 2096 19771
rect 2044 19728 2096 19737
rect 4344 19728 4396 19780
rect 5080 19796 5132 19848
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 6828 19728 6880 19780
rect 7380 19796 7432 19848
rect 7656 19839 7708 19848
rect 7656 19805 7665 19839
rect 7665 19805 7699 19839
rect 7699 19805 7708 19839
rect 7656 19796 7708 19805
rect 5448 19660 5500 19712
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 7288 19660 7340 19712
rect 8668 19796 8720 19848
rect 8760 19796 8812 19848
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 11888 19864 11940 19916
rect 12532 19864 12584 19916
rect 15108 19907 15160 19916
rect 15108 19873 15117 19907
rect 15117 19873 15151 19907
rect 15151 19873 15160 19907
rect 15108 19864 15160 19873
rect 16304 20000 16356 20052
rect 16120 19932 16172 19984
rect 17500 20000 17552 20052
rect 18328 20000 18380 20052
rect 8944 19660 8996 19712
rect 9036 19660 9088 19712
rect 11336 19796 11388 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 12808 19728 12860 19780
rect 15384 19796 15436 19848
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16304 19864 16356 19916
rect 18880 19975 18932 19984
rect 18880 19941 18889 19975
rect 18889 19941 18923 19975
rect 18923 19941 18932 19975
rect 18880 19932 18932 19941
rect 20628 19932 20680 19984
rect 25964 19932 26016 19984
rect 16120 19796 16172 19805
rect 13360 19660 13412 19712
rect 15384 19660 15436 19712
rect 16028 19660 16080 19712
rect 16580 19771 16632 19780
rect 16580 19737 16589 19771
rect 16589 19737 16623 19771
rect 16623 19737 16632 19771
rect 16580 19728 16632 19737
rect 19340 19864 19392 19916
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 24124 19907 24176 19916
rect 24124 19873 24133 19907
rect 24133 19873 24167 19907
rect 24167 19873 24176 19907
rect 24124 19864 24176 19873
rect 24676 19864 24728 19916
rect 24860 19796 24912 19848
rect 26056 19796 26108 19848
rect 23848 19771 23900 19780
rect 23848 19737 23857 19771
rect 23857 19737 23891 19771
rect 23891 19737 23900 19771
rect 23848 19728 23900 19737
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 19616 19660 19668 19712
rect 19800 19703 19852 19712
rect 19800 19669 19809 19703
rect 19809 19669 19843 19703
rect 19843 19669 19852 19703
rect 19800 19660 19852 19669
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 21548 19660 21600 19712
rect 23112 19660 23164 19712
rect 24400 19703 24452 19712
rect 24400 19669 24409 19703
rect 24409 19669 24443 19703
rect 24443 19669 24452 19703
rect 24400 19660 24452 19669
rect 25228 19660 25280 19712
rect 4703 19558 4755 19610
rect 4767 19558 4819 19610
rect 4831 19558 4883 19610
rect 4895 19558 4947 19610
rect 4959 19558 5011 19610
rect 10890 19558 10942 19610
rect 10954 19558 11006 19610
rect 11018 19558 11070 19610
rect 11082 19558 11134 19610
rect 11146 19558 11198 19610
rect 17077 19558 17129 19610
rect 17141 19558 17193 19610
rect 17205 19558 17257 19610
rect 17269 19558 17321 19610
rect 17333 19558 17385 19610
rect 23264 19558 23316 19610
rect 23328 19558 23380 19610
rect 23392 19558 23444 19610
rect 23456 19558 23508 19610
rect 23520 19558 23572 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2044 19456 2096 19508
rect 2596 19456 2648 19508
rect 2688 19456 2740 19508
rect 1492 19363 1544 19372
rect 1492 19329 1501 19363
rect 1501 19329 1535 19363
rect 1535 19329 1544 19363
rect 1492 19320 1544 19329
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 3516 19388 3568 19440
rect 4344 19456 4396 19508
rect 4436 19388 4488 19440
rect 4528 19388 4580 19440
rect 3608 19252 3660 19304
rect 1860 19184 1912 19236
rect 2136 19159 2188 19168
rect 2136 19125 2145 19159
rect 2145 19125 2179 19159
rect 2179 19125 2188 19159
rect 2136 19116 2188 19125
rect 4804 19320 4856 19372
rect 4528 19252 4580 19304
rect 4620 19184 4672 19236
rect 6460 19456 6512 19508
rect 7656 19456 7708 19508
rect 8300 19456 8352 19508
rect 10692 19456 10744 19508
rect 13084 19456 13136 19508
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 5908 19388 5960 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 7196 19388 7248 19440
rect 8576 19388 8628 19440
rect 12716 19388 12768 19440
rect 14832 19388 14884 19440
rect 15568 19388 15620 19440
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 6920 19320 6972 19372
rect 7104 19320 7156 19372
rect 7564 19320 7616 19372
rect 8392 19252 8444 19304
rect 8484 19252 8536 19304
rect 9128 19252 9180 19304
rect 16580 19388 16632 19440
rect 17040 19388 17092 19440
rect 12348 19252 12400 19304
rect 11612 19184 11664 19236
rect 12624 19295 12676 19304
rect 12624 19261 12633 19295
rect 12633 19261 12667 19295
rect 12667 19261 12676 19295
rect 12624 19252 12676 19261
rect 12992 19320 13044 19372
rect 14188 19320 14240 19372
rect 15384 19320 15436 19372
rect 16120 19320 16172 19372
rect 16304 19363 16356 19372
rect 16304 19329 16313 19363
rect 16313 19329 16347 19363
rect 16347 19329 16356 19363
rect 16304 19320 16356 19329
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 4528 19116 4580 19168
rect 5172 19116 5224 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 9772 19116 9824 19168
rect 9956 19116 10008 19168
rect 10692 19116 10744 19168
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 12808 19184 12860 19236
rect 14372 19252 14424 19304
rect 15108 19252 15160 19304
rect 15200 19252 15252 19304
rect 15660 19252 15712 19304
rect 15936 19252 15988 19304
rect 18052 19431 18104 19440
rect 18052 19397 18061 19431
rect 18061 19397 18095 19431
rect 18095 19397 18104 19431
rect 18052 19388 18104 19397
rect 19340 19388 19392 19440
rect 18512 19252 18564 19304
rect 19800 19456 19852 19508
rect 19892 19456 19944 19508
rect 23112 19456 23164 19508
rect 25228 19499 25280 19508
rect 25228 19465 25237 19499
rect 25237 19465 25271 19499
rect 25271 19465 25280 19499
rect 25228 19456 25280 19465
rect 22192 19431 22244 19440
rect 22192 19397 22201 19431
rect 22201 19397 22235 19431
rect 22235 19397 22244 19431
rect 22192 19388 22244 19397
rect 21640 19363 21692 19372
rect 21640 19329 21649 19363
rect 21649 19329 21683 19363
rect 21683 19329 21692 19363
rect 21640 19320 21692 19329
rect 23664 19388 23716 19440
rect 24400 19388 24452 19440
rect 14740 19184 14792 19236
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 14924 19116 14976 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 15844 19227 15896 19236
rect 15844 19193 15853 19227
rect 15853 19193 15887 19227
rect 15887 19193 15896 19227
rect 15844 19184 15896 19193
rect 16672 19116 16724 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 19432 19116 19484 19168
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 23020 19252 23072 19304
rect 25780 19320 25832 19372
rect 21180 19184 21232 19236
rect 23480 19184 23532 19236
rect 20536 19116 20588 19168
rect 23112 19116 23164 19168
rect 4043 19014 4095 19066
rect 4107 19014 4159 19066
rect 4171 19014 4223 19066
rect 4235 19014 4287 19066
rect 4299 19014 4351 19066
rect 10230 19014 10282 19066
rect 10294 19014 10346 19066
rect 10358 19014 10410 19066
rect 10422 19014 10474 19066
rect 10486 19014 10538 19066
rect 16417 19014 16469 19066
rect 16481 19014 16533 19066
rect 16545 19014 16597 19066
rect 16609 19014 16661 19066
rect 16673 19014 16725 19066
rect 22604 19014 22656 19066
rect 22668 19014 22720 19066
rect 22732 19014 22784 19066
rect 22796 19014 22848 19066
rect 22860 19014 22912 19066
rect 3792 18955 3844 18964
rect 3792 18921 3801 18955
rect 3801 18921 3835 18955
rect 3835 18921 3844 18955
rect 3792 18912 3844 18921
rect 4344 18912 4396 18964
rect 4896 18912 4948 18964
rect 5080 18912 5132 18964
rect 5356 18912 5408 18964
rect 6644 18912 6696 18964
rect 8024 18912 8076 18964
rect 4252 18844 4304 18896
rect 3608 18776 3660 18828
rect 4344 18819 4396 18828
rect 4344 18785 4353 18819
rect 4353 18785 4387 18819
rect 4387 18785 4396 18819
rect 4344 18776 4396 18785
rect 5264 18844 5316 18896
rect 5816 18844 5868 18896
rect 7380 18844 7432 18896
rect 7656 18844 7708 18896
rect 9496 18912 9548 18964
rect 9772 18912 9824 18964
rect 11612 18955 11664 18964
rect 11612 18921 11621 18955
rect 11621 18921 11655 18955
rect 11655 18921 11664 18955
rect 11612 18912 11664 18921
rect 14188 18955 14240 18964
rect 14188 18921 14197 18955
rect 14197 18921 14231 18955
rect 14231 18921 14240 18955
rect 14188 18912 14240 18921
rect 14464 18912 14516 18964
rect 14740 18912 14792 18964
rect 15292 18912 15344 18964
rect 15844 18955 15896 18964
rect 15844 18921 15853 18955
rect 15853 18921 15887 18955
rect 15887 18921 15896 18955
rect 15844 18912 15896 18921
rect 15936 18912 15988 18964
rect 8300 18887 8352 18896
rect 8300 18853 8309 18887
rect 8309 18853 8343 18887
rect 8343 18853 8352 18887
rect 8300 18844 8352 18853
rect 8668 18844 8720 18896
rect 4620 18708 4672 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 7840 18776 7892 18828
rect 8484 18776 8536 18828
rect 9036 18776 9088 18828
rect 5724 18708 5776 18760
rect 6092 18708 6144 18760
rect 6920 18708 6972 18760
rect 7564 18708 7616 18760
rect 11336 18776 11388 18828
rect 15476 18844 15528 18896
rect 15844 18819 15896 18828
rect 15844 18785 15850 18819
rect 15850 18785 15884 18819
rect 15884 18785 15896 18819
rect 15844 18776 15896 18785
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 13912 18708 13964 18760
rect 4160 18683 4212 18692
rect 4160 18649 4169 18683
rect 4169 18649 4203 18683
rect 4203 18649 4212 18683
rect 4160 18640 4212 18649
rect 5356 18640 5408 18692
rect 9036 18640 9088 18692
rect 10140 18683 10192 18692
rect 10140 18649 10149 18683
rect 10149 18649 10183 18683
rect 10183 18649 10192 18683
rect 10140 18640 10192 18649
rect 10600 18640 10652 18692
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 4620 18572 4672 18624
rect 4896 18572 4948 18624
rect 14740 18640 14792 18692
rect 11796 18615 11848 18624
rect 11796 18581 11805 18615
rect 11805 18581 11839 18615
rect 11839 18581 11848 18615
rect 11796 18572 11848 18581
rect 11980 18572 12032 18624
rect 15108 18708 15160 18760
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 15568 18708 15620 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16304 18912 16356 18964
rect 18236 18912 18288 18964
rect 19340 18912 19392 18964
rect 19892 18912 19944 18964
rect 19984 18912 20036 18964
rect 24492 18912 24544 18964
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 25412 18955 25464 18964
rect 25412 18921 25421 18955
rect 25421 18921 25455 18955
rect 25455 18921 25464 18955
rect 25412 18912 25464 18921
rect 14924 18640 14976 18692
rect 15384 18640 15436 18692
rect 16488 18708 16540 18760
rect 16672 18708 16724 18760
rect 16764 18708 16816 18760
rect 17500 18708 17552 18760
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 18788 18819 18840 18828
rect 18788 18785 18797 18819
rect 18797 18785 18831 18819
rect 18831 18785 18840 18819
rect 18788 18776 18840 18785
rect 23940 18844 23992 18896
rect 19340 18776 19392 18828
rect 19616 18776 19668 18828
rect 20536 18776 20588 18828
rect 15108 18572 15160 18624
rect 16856 18640 16908 18692
rect 17776 18640 17828 18692
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 23480 18776 23532 18828
rect 23664 18776 23716 18828
rect 23020 18708 23072 18760
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 25228 18751 25280 18760
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 19892 18640 19944 18692
rect 21180 18640 21232 18692
rect 21548 18640 21600 18692
rect 17040 18572 17092 18624
rect 17592 18572 17644 18624
rect 22284 18572 22336 18624
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 4703 18470 4755 18522
rect 4767 18470 4819 18522
rect 4831 18470 4883 18522
rect 4895 18470 4947 18522
rect 4959 18470 5011 18522
rect 10890 18470 10942 18522
rect 10954 18470 11006 18522
rect 11018 18470 11070 18522
rect 11082 18470 11134 18522
rect 11146 18470 11198 18522
rect 17077 18470 17129 18522
rect 17141 18470 17193 18522
rect 17205 18470 17257 18522
rect 17269 18470 17321 18522
rect 17333 18470 17385 18522
rect 23264 18470 23316 18522
rect 23328 18470 23380 18522
rect 23392 18470 23444 18522
rect 23456 18470 23508 18522
rect 23520 18470 23572 18522
rect 4528 18368 4580 18420
rect 6368 18300 6420 18352
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 3056 18232 3108 18284
rect 7012 18275 7064 18284
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 2228 18096 2280 18148
rect 7196 18164 7248 18216
rect 8944 18411 8996 18420
rect 8944 18377 8953 18411
rect 8953 18377 8987 18411
rect 8987 18377 8996 18411
rect 8944 18368 8996 18377
rect 9220 18368 9272 18420
rect 10140 18368 10192 18420
rect 10692 18368 10744 18420
rect 12808 18368 12860 18420
rect 13912 18368 13964 18420
rect 15752 18368 15804 18420
rect 15936 18368 15988 18420
rect 16488 18368 16540 18420
rect 16672 18368 16724 18420
rect 19984 18368 20036 18420
rect 20996 18368 21048 18420
rect 21640 18368 21692 18420
rect 22284 18411 22336 18420
rect 22284 18377 22293 18411
rect 22293 18377 22327 18411
rect 22327 18377 22336 18411
rect 22284 18368 22336 18377
rect 23112 18368 23164 18420
rect 7564 18232 7616 18284
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 8668 18232 8720 18284
rect 12440 18300 12492 18352
rect 14648 18300 14700 18352
rect 15384 18343 15436 18352
rect 15384 18309 15393 18343
rect 15393 18309 15427 18343
rect 15427 18309 15436 18343
rect 15384 18300 15436 18309
rect 15476 18300 15528 18352
rect 15844 18300 15896 18352
rect 16396 18300 16448 18352
rect 17408 18300 17460 18352
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2044 18028 2096 18080
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 6092 18028 6144 18037
rect 7104 18071 7156 18080
rect 7104 18037 7113 18071
rect 7113 18037 7147 18071
rect 7147 18037 7156 18071
rect 7104 18028 7156 18037
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 11336 18164 11388 18216
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15108 18232 15160 18284
rect 15200 18232 15252 18284
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 17040 18232 17092 18284
rect 17500 18232 17552 18284
rect 17776 18232 17828 18284
rect 19340 18232 19392 18284
rect 20536 18232 20588 18284
rect 23296 18300 23348 18352
rect 24952 18300 25004 18352
rect 25964 18300 26016 18352
rect 7932 18028 7984 18080
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 15384 18028 15436 18080
rect 16764 18207 16816 18216
rect 16764 18173 16773 18207
rect 16773 18173 16807 18207
rect 16807 18173 16816 18207
rect 16764 18164 16816 18173
rect 15844 18096 15896 18148
rect 17776 18096 17828 18148
rect 21640 18096 21692 18148
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 17040 18028 17092 18037
rect 17132 18028 17184 18080
rect 17316 18071 17368 18080
rect 17316 18037 17325 18071
rect 17325 18037 17359 18071
rect 17359 18037 17368 18071
rect 17316 18028 17368 18037
rect 18512 18028 18564 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 22376 18207 22428 18216
rect 22376 18173 22385 18207
rect 22385 18173 22419 18207
rect 22419 18173 22428 18207
rect 22376 18164 22428 18173
rect 23020 18164 23072 18216
rect 24492 18028 24544 18080
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 25320 18071 25372 18080
rect 25320 18037 25329 18071
rect 25329 18037 25363 18071
rect 25363 18037 25372 18071
rect 25320 18028 25372 18037
rect 4043 17926 4095 17978
rect 4107 17926 4159 17978
rect 4171 17926 4223 17978
rect 4235 17926 4287 17978
rect 4299 17926 4351 17978
rect 10230 17926 10282 17978
rect 10294 17926 10346 17978
rect 10358 17926 10410 17978
rect 10422 17926 10474 17978
rect 10486 17926 10538 17978
rect 16417 17926 16469 17978
rect 16481 17926 16533 17978
rect 16545 17926 16597 17978
rect 16609 17926 16661 17978
rect 16673 17926 16725 17978
rect 22604 17926 22656 17978
rect 22668 17926 22720 17978
rect 22732 17926 22784 17978
rect 22796 17926 22848 17978
rect 22860 17926 22912 17978
rect 4436 17824 4488 17876
rect 6920 17824 6972 17876
rect 7380 17824 7432 17876
rect 7564 17824 7616 17876
rect 8116 17824 8168 17876
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 1676 17688 1728 17697
rect 2044 17688 2096 17740
rect 3700 17688 3752 17740
rect 9036 17867 9088 17876
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 13268 17824 13320 17876
rect 13912 17824 13964 17876
rect 15568 17824 15620 17876
rect 7932 17688 7984 17740
rect 4068 17620 4120 17672
rect 2228 17552 2280 17604
rect 5264 17663 5316 17672
rect 5264 17629 5273 17663
rect 5273 17629 5307 17663
rect 5307 17629 5316 17663
rect 5264 17620 5316 17629
rect 7012 17620 7064 17672
rect 7380 17663 7432 17672
rect 7380 17629 7389 17663
rect 7389 17629 7423 17663
rect 7423 17629 7432 17663
rect 7380 17620 7432 17629
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 2872 17484 2924 17536
rect 3976 17484 4028 17536
rect 7104 17484 7156 17536
rect 8300 17620 8352 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 9036 17620 9088 17672
rect 9680 17688 9732 17740
rect 14740 17688 14792 17740
rect 14832 17688 14884 17740
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 15476 17688 15528 17740
rect 9496 17595 9548 17604
rect 9496 17561 9505 17595
rect 9505 17561 9539 17595
rect 9539 17561 9548 17595
rect 9496 17552 9548 17561
rect 9680 17552 9732 17604
rect 11704 17595 11756 17604
rect 11704 17561 11713 17595
rect 11713 17561 11747 17595
rect 11747 17561 11756 17595
rect 11704 17552 11756 17561
rect 7932 17484 7984 17536
rect 8392 17484 8444 17536
rect 13728 17484 13780 17536
rect 14464 17552 14516 17604
rect 15384 17552 15436 17604
rect 15936 17824 15988 17876
rect 19432 17824 19484 17876
rect 19616 17824 19668 17876
rect 17316 17756 17368 17808
rect 22468 17824 22520 17876
rect 23204 17824 23256 17876
rect 25136 17824 25188 17876
rect 19892 17731 19944 17740
rect 19892 17697 19901 17731
rect 19901 17697 19935 17731
rect 19935 17697 19944 17731
rect 19892 17688 19944 17697
rect 22192 17688 22244 17740
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16304 17620 16356 17672
rect 17040 17620 17092 17672
rect 20536 17663 20588 17672
rect 20536 17629 20545 17663
rect 20545 17629 20579 17663
rect 20579 17629 20588 17663
rect 20536 17620 20588 17629
rect 23940 17799 23992 17808
rect 23940 17765 23949 17799
rect 23949 17765 23983 17799
rect 23983 17765 23992 17799
rect 23940 17756 23992 17765
rect 24400 17799 24452 17808
rect 24400 17765 24409 17799
rect 24409 17765 24443 17799
rect 24443 17765 24452 17799
rect 24400 17756 24452 17765
rect 24676 17756 24728 17808
rect 19800 17552 19852 17604
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 21272 17552 21324 17604
rect 16028 17484 16080 17536
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 21824 17484 21876 17536
rect 22836 17552 22888 17604
rect 23664 17731 23716 17740
rect 23664 17697 23673 17731
rect 23673 17697 23707 17731
rect 23707 17697 23716 17731
rect 23664 17688 23716 17697
rect 24124 17688 24176 17740
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 23296 17620 23348 17672
rect 24032 17620 24084 17672
rect 22652 17484 22704 17536
rect 25136 17484 25188 17536
rect 4703 17382 4755 17434
rect 4767 17382 4819 17434
rect 4831 17382 4883 17434
rect 4895 17382 4947 17434
rect 4959 17382 5011 17434
rect 10890 17382 10942 17434
rect 10954 17382 11006 17434
rect 11018 17382 11070 17434
rect 11082 17382 11134 17434
rect 11146 17382 11198 17434
rect 17077 17382 17129 17434
rect 17141 17382 17193 17434
rect 17205 17382 17257 17434
rect 17269 17382 17321 17434
rect 17333 17382 17385 17434
rect 23264 17382 23316 17434
rect 23328 17382 23380 17434
rect 23392 17382 23444 17434
rect 23456 17382 23508 17434
rect 23520 17382 23572 17434
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 2872 17280 2924 17332
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3700 17280 3752 17332
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 940 17076 992 17128
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 2780 17144 2832 17196
rect 3148 17119 3200 17128
rect 3148 17085 3157 17119
rect 3157 17085 3191 17119
rect 3191 17085 3200 17119
rect 3148 17076 3200 17085
rect 4436 17280 4488 17332
rect 5908 17280 5960 17332
rect 8576 17280 8628 17332
rect 8760 17280 8812 17332
rect 12440 17280 12492 17332
rect 14740 17280 14792 17332
rect 15660 17280 15712 17332
rect 16212 17280 16264 17332
rect 20812 17280 20864 17332
rect 22652 17280 22704 17332
rect 22836 17280 22888 17332
rect 23112 17280 23164 17332
rect 4068 17144 4120 17196
rect 4620 17255 4672 17264
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 4620 17212 4672 17221
rect 6000 17212 6052 17264
rect 7196 17212 7248 17264
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 1860 16983 1912 16992
rect 1860 16949 1869 16983
rect 1869 16949 1903 16983
rect 1903 16949 1912 16983
rect 1860 16940 1912 16949
rect 2044 16940 2096 16992
rect 3516 17051 3568 17060
rect 3516 17017 3525 17051
rect 3525 17017 3559 17051
rect 3559 17017 3568 17051
rect 3516 17008 3568 17017
rect 3700 17008 3752 17060
rect 3976 16940 4028 16992
rect 5724 17008 5776 17060
rect 6092 16940 6144 16992
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 7656 17187 7708 17196
rect 7656 17153 7665 17187
rect 7665 17153 7699 17187
rect 7699 17153 7708 17187
rect 7656 17144 7708 17153
rect 8024 17144 8076 17196
rect 8392 17255 8444 17264
rect 8392 17221 8401 17255
rect 8401 17221 8435 17255
rect 8435 17221 8444 17255
rect 8392 17212 8444 17221
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 12808 17212 12860 17264
rect 15568 17212 15620 17264
rect 15844 17212 15896 17264
rect 16028 17212 16080 17264
rect 7932 17076 7984 17128
rect 8576 17008 8628 17060
rect 9588 17008 9640 17060
rect 12072 17119 12124 17128
rect 12072 17085 12081 17119
rect 12081 17085 12115 17119
rect 12115 17085 12124 17119
rect 12072 17076 12124 17085
rect 12624 17144 12676 17196
rect 13820 17076 13872 17128
rect 8392 16940 8444 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 15752 17144 15804 17196
rect 19156 17144 19208 17196
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 20352 17144 20404 17196
rect 15292 17076 15344 17128
rect 16856 17076 16908 17128
rect 21180 17076 21232 17128
rect 21640 17076 21692 17128
rect 20628 17008 20680 17060
rect 12440 16940 12492 16992
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 15568 16940 15620 16992
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 18696 16940 18748 16992
rect 19616 16983 19668 16992
rect 19616 16949 19625 16983
rect 19625 16949 19659 16983
rect 19659 16949 19668 16983
rect 19616 16940 19668 16949
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 22376 17119 22428 17128
rect 22376 17085 22385 17119
rect 22385 17085 22419 17119
rect 22419 17085 22428 17119
rect 22376 17076 22428 17085
rect 24400 17280 24452 17332
rect 23664 17212 23716 17264
rect 23940 17008 23992 17060
rect 24584 17008 24636 17060
rect 25688 17076 25740 17128
rect 25964 17008 26016 17060
rect 24032 16940 24084 16992
rect 24860 16940 24912 16992
rect 4043 16838 4095 16890
rect 4107 16838 4159 16890
rect 4171 16838 4223 16890
rect 4235 16838 4287 16890
rect 4299 16838 4351 16890
rect 10230 16838 10282 16890
rect 10294 16838 10346 16890
rect 10358 16838 10410 16890
rect 10422 16838 10474 16890
rect 10486 16838 10538 16890
rect 16417 16838 16469 16890
rect 16481 16838 16533 16890
rect 16545 16838 16597 16890
rect 16609 16838 16661 16890
rect 16673 16838 16725 16890
rect 22604 16838 22656 16890
rect 22668 16838 22720 16890
rect 22732 16838 22784 16890
rect 22796 16838 22848 16890
rect 22860 16838 22912 16890
rect 1676 16736 1728 16788
rect 2872 16736 2924 16788
rect 3516 16736 3568 16788
rect 4252 16668 4304 16720
rect 4528 16711 4580 16720
rect 4528 16677 4537 16711
rect 4537 16677 4571 16711
rect 4571 16677 4580 16711
rect 4528 16668 4580 16677
rect 6000 16779 6052 16788
rect 6000 16745 6009 16779
rect 6009 16745 6043 16779
rect 6043 16745 6052 16779
rect 6000 16736 6052 16745
rect 6368 16779 6420 16788
rect 6368 16745 6377 16779
rect 6377 16745 6411 16779
rect 6411 16745 6420 16779
rect 6368 16736 6420 16745
rect 11060 16736 11112 16788
rect 11152 16736 11204 16788
rect 5540 16668 5592 16720
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 3700 16532 3752 16584
rect 5448 16600 5500 16652
rect 3792 16464 3844 16516
rect 4620 16464 4672 16516
rect 4068 16396 4120 16448
rect 5448 16507 5500 16516
rect 5448 16473 5457 16507
rect 5457 16473 5491 16507
rect 5491 16473 5500 16507
rect 5448 16464 5500 16473
rect 9588 16600 9640 16652
rect 10600 16668 10652 16720
rect 10416 16600 10468 16652
rect 12072 16600 12124 16652
rect 16948 16736 17000 16788
rect 14556 16668 14608 16720
rect 16856 16668 16908 16720
rect 14924 16600 14976 16652
rect 15568 16600 15620 16652
rect 15752 16600 15804 16652
rect 8024 16464 8076 16516
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 8760 16575 8812 16584
rect 8760 16541 8769 16575
rect 8769 16541 8803 16575
rect 8803 16541 8812 16575
rect 8760 16532 8812 16541
rect 8944 16532 8996 16584
rect 10692 16464 10744 16516
rect 12440 16532 12492 16584
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 11336 16464 11388 16516
rect 13452 16464 13504 16516
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 19800 16736 19852 16788
rect 20904 16736 20956 16788
rect 18236 16643 18288 16652
rect 18236 16609 18245 16643
rect 18245 16609 18279 16643
rect 18279 16609 18288 16643
rect 18236 16600 18288 16609
rect 18696 16600 18748 16652
rect 20628 16643 20680 16652
rect 20628 16609 20637 16643
rect 20637 16609 20671 16643
rect 20671 16609 20680 16643
rect 20628 16600 20680 16609
rect 18144 16532 18196 16584
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 19800 16532 19852 16584
rect 20352 16532 20404 16584
rect 21916 16736 21968 16788
rect 22192 16668 22244 16720
rect 22376 16668 22428 16720
rect 23664 16668 23716 16720
rect 24676 16668 24728 16720
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 10048 16396 10100 16448
rect 12624 16396 12676 16448
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 14188 16396 14240 16448
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15384 16464 15436 16516
rect 17776 16396 17828 16448
rect 19432 16464 19484 16516
rect 21824 16532 21876 16584
rect 23848 16600 23900 16652
rect 24952 16600 25004 16652
rect 19064 16396 19116 16448
rect 20904 16396 20956 16448
rect 22284 16464 22336 16516
rect 21180 16396 21232 16448
rect 22008 16396 22060 16448
rect 23940 16532 23992 16584
rect 22836 16464 22888 16516
rect 24860 16532 24912 16584
rect 22468 16396 22520 16448
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 25228 16396 25280 16448
rect 4703 16294 4755 16346
rect 4767 16294 4819 16346
rect 4831 16294 4883 16346
rect 4895 16294 4947 16346
rect 4959 16294 5011 16346
rect 10890 16294 10942 16346
rect 10954 16294 11006 16346
rect 11018 16294 11070 16346
rect 11082 16294 11134 16346
rect 11146 16294 11198 16346
rect 17077 16294 17129 16346
rect 17141 16294 17193 16346
rect 17205 16294 17257 16346
rect 17269 16294 17321 16346
rect 17333 16294 17385 16346
rect 23264 16294 23316 16346
rect 23328 16294 23380 16346
rect 23392 16294 23444 16346
rect 23456 16294 23508 16346
rect 23520 16294 23572 16346
rect 3608 16192 3660 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 4528 16192 4580 16244
rect 7840 16192 7892 16244
rect 8024 16192 8076 16244
rect 8576 16192 8628 16244
rect 9220 16192 9272 16244
rect 9496 16192 9548 16244
rect 10784 16192 10836 16244
rect 10968 16192 11020 16244
rect 2780 16124 2832 16176
rect 4068 16124 4120 16176
rect 4620 16124 4672 16176
rect 11704 16192 11756 16244
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 940 15852 992 15904
rect 2504 15988 2556 16040
rect 2872 15963 2924 15972
rect 2872 15929 2881 15963
rect 2881 15929 2915 15963
rect 2915 15929 2924 15963
rect 2872 15920 2924 15929
rect 3056 15988 3108 16040
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 6920 16056 6972 16108
rect 9312 16056 9364 16108
rect 11428 16124 11480 16176
rect 11520 16124 11572 16176
rect 11888 16124 11940 16176
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 11060 16056 11112 16108
rect 11796 16099 11848 16108
rect 11796 16065 11805 16099
rect 11805 16065 11839 16099
rect 11839 16065 11848 16099
rect 11796 16056 11848 16065
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 12624 16124 12676 16176
rect 15476 16124 15528 16176
rect 17500 16192 17552 16244
rect 17776 16192 17828 16244
rect 16212 16124 16264 16176
rect 17592 16124 17644 16176
rect 18236 16124 18288 16176
rect 18972 16235 19024 16244
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 20352 16192 20404 16244
rect 22008 16192 22060 16244
rect 3148 15920 3200 15972
rect 10416 15988 10468 16040
rect 10600 15920 10652 15972
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 11336 15988 11388 16040
rect 11152 15963 11204 15972
rect 11152 15929 11161 15963
rect 11161 15929 11195 15963
rect 11195 15929 11204 15963
rect 11152 15920 11204 15929
rect 12716 16031 12768 16040
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 12716 15988 12768 15997
rect 12808 15988 12860 16040
rect 19340 16056 19392 16108
rect 19616 16056 19668 16108
rect 19800 16056 19852 16108
rect 21824 16167 21876 16176
rect 21824 16133 21833 16167
rect 21833 16133 21867 16167
rect 21867 16133 21876 16167
rect 21824 16124 21876 16133
rect 15292 15988 15344 16040
rect 15752 15988 15804 16040
rect 5632 15852 5684 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 10048 15852 10100 15904
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 17592 15988 17644 16040
rect 18144 15988 18196 16040
rect 18788 15988 18840 16040
rect 21088 15988 21140 16040
rect 18512 15920 18564 15972
rect 19616 15920 19668 15972
rect 13452 15852 13504 15904
rect 14188 15895 14240 15904
rect 14188 15861 14197 15895
rect 14197 15861 14231 15895
rect 14231 15861 14240 15895
rect 14188 15852 14240 15861
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 15936 15852 15988 15904
rect 16212 15852 16264 15904
rect 19340 15852 19392 15904
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 19892 15852 19944 15904
rect 20720 15852 20772 15904
rect 21916 16056 21968 16108
rect 22836 16235 22888 16244
rect 22836 16201 22845 16235
rect 22845 16201 22879 16235
rect 22879 16201 22888 16235
rect 22836 16192 22888 16201
rect 23388 16192 23440 16244
rect 23848 16192 23900 16244
rect 25228 16124 25280 16176
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 22100 15988 22152 16040
rect 23388 16031 23440 16040
rect 23388 15997 23397 16031
rect 23397 15997 23431 16031
rect 23431 15997 23440 16031
rect 23388 15988 23440 15997
rect 22192 15963 22244 15972
rect 22192 15929 22201 15963
rect 22201 15929 22235 15963
rect 22235 15929 22244 15963
rect 22192 15920 22244 15929
rect 22284 15920 22336 15972
rect 23020 15920 23072 15972
rect 25228 15988 25280 16040
rect 26148 16192 26200 16244
rect 25504 15852 25556 15904
rect 4043 15750 4095 15802
rect 4107 15750 4159 15802
rect 4171 15750 4223 15802
rect 4235 15750 4287 15802
rect 4299 15750 4351 15802
rect 10230 15750 10282 15802
rect 10294 15750 10346 15802
rect 10358 15750 10410 15802
rect 10422 15750 10474 15802
rect 10486 15750 10538 15802
rect 16417 15750 16469 15802
rect 16481 15750 16533 15802
rect 16545 15750 16597 15802
rect 16609 15750 16661 15802
rect 16673 15750 16725 15802
rect 22604 15750 22656 15802
rect 22668 15750 22720 15802
rect 22732 15750 22784 15802
rect 22796 15750 22848 15802
rect 22860 15750 22912 15802
rect 2044 15444 2096 15496
rect 3792 15580 3844 15632
rect 3516 15512 3568 15564
rect 6920 15648 6972 15700
rect 9312 15648 9364 15700
rect 9588 15648 9640 15700
rect 9956 15648 10008 15700
rect 10876 15648 10928 15700
rect 12624 15648 12676 15700
rect 12716 15648 12768 15700
rect 7932 15580 7984 15632
rect 19064 15648 19116 15700
rect 19892 15648 19944 15700
rect 20904 15648 20956 15700
rect 22192 15648 22244 15700
rect 17500 15580 17552 15632
rect 18880 15623 18932 15632
rect 18880 15589 18889 15623
rect 18889 15589 18923 15623
rect 18923 15589 18932 15623
rect 18880 15580 18932 15589
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 3332 15444 3384 15496
rect 5632 15512 5684 15564
rect 11244 15512 11296 15564
rect 11336 15512 11388 15564
rect 8208 15487 8260 15496
rect 2780 15308 2832 15360
rect 3516 15308 3568 15360
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 9128 15444 9180 15496
rect 9956 15444 10008 15496
rect 10968 15444 11020 15496
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11612 15444 11664 15496
rect 13176 15512 13228 15564
rect 14556 15512 14608 15564
rect 15292 15512 15344 15564
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 5724 15376 5776 15428
rect 16120 15376 16172 15428
rect 16304 15376 16356 15428
rect 17592 15376 17644 15428
rect 7012 15308 7064 15360
rect 10048 15308 10100 15360
rect 11152 15308 11204 15360
rect 15384 15308 15436 15360
rect 16948 15308 17000 15360
rect 18788 15376 18840 15428
rect 19800 15376 19852 15428
rect 22284 15512 22336 15564
rect 23388 15648 23440 15700
rect 23940 15648 23992 15700
rect 25412 15691 25464 15700
rect 25412 15657 25421 15691
rect 25421 15657 25455 15691
rect 25455 15657 25464 15691
rect 25412 15648 25464 15657
rect 23756 15512 23808 15564
rect 23940 15512 23992 15564
rect 24400 15512 24452 15564
rect 24492 15444 24544 15496
rect 26240 15444 26292 15496
rect 22284 15376 22336 15428
rect 22468 15376 22520 15428
rect 18880 15308 18932 15360
rect 22008 15308 22060 15360
rect 24216 15351 24268 15360
rect 24216 15317 24225 15351
rect 24225 15317 24259 15351
rect 24259 15317 24268 15351
rect 24216 15308 24268 15317
rect 4703 15206 4755 15258
rect 4767 15206 4819 15258
rect 4831 15206 4883 15258
rect 4895 15206 4947 15258
rect 4959 15206 5011 15258
rect 10890 15206 10942 15258
rect 10954 15206 11006 15258
rect 11018 15206 11070 15258
rect 11082 15206 11134 15258
rect 11146 15206 11198 15258
rect 17077 15206 17129 15258
rect 17141 15206 17193 15258
rect 17205 15206 17257 15258
rect 17269 15206 17321 15258
rect 17333 15206 17385 15258
rect 23264 15206 23316 15258
rect 23328 15206 23380 15258
rect 23392 15206 23444 15258
rect 23456 15206 23508 15258
rect 23520 15206 23572 15258
rect 1676 15104 1728 15156
rect 2780 15104 2832 15156
rect 5908 15104 5960 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 3516 15036 3568 15088
rect 3884 15036 3936 15088
rect 2964 14968 3016 15020
rect 3148 14968 3200 15020
rect 5448 14968 5500 15020
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 2412 14764 2464 14816
rect 3332 14875 3384 14884
rect 3332 14841 3341 14875
rect 3341 14841 3375 14875
rect 3375 14841 3384 14875
rect 3332 14832 3384 14841
rect 5540 14875 5592 14884
rect 5540 14841 5549 14875
rect 5549 14841 5583 14875
rect 5583 14841 5592 14875
rect 5540 14832 5592 14841
rect 7656 14968 7708 15020
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 8484 14900 8536 14952
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5080 14764 5132 14816
rect 5632 14764 5684 14816
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 10784 14900 10836 14909
rect 10692 14832 10744 14884
rect 11060 14875 11112 14884
rect 11060 14841 11069 14875
rect 11069 14841 11103 14875
rect 11103 14841 11112 14875
rect 11060 14832 11112 14841
rect 11244 14764 11296 14816
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 13544 14832 13596 14884
rect 17408 15104 17460 15156
rect 18236 15147 18288 15156
rect 18236 15113 18245 15147
rect 18245 15113 18279 15147
rect 18279 15113 18288 15147
rect 18236 15104 18288 15113
rect 19156 15147 19208 15156
rect 19156 15113 19165 15147
rect 19165 15113 19199 15147
rect 19199 15113 19208 15147
rect 19156 15104 19208 15113
rect 19800 15147 19852 15156
rect 19800 15113 19809 15147
rect 19809 15113 19843 15147
rect 19843 15113 19852 15147
rect 19800 15104 19852 15113
rect 20720 15104 20772 15156
rect 22376 15147 22428 15156
rect 22376 15113 22385 15147
rect 22385 15113 22419 15147
rect 22419 15113 22428 15147
rect 22376 15104 22428 15113
rect 24216 15104 24268 15156
rect 24952 15104 25004 15156
rect 15016 15036 15068 15088
rect 15200 15036 15252 15088
rect 16212 15036 16264 15088
rect 15384 15011 15436 15020
rect 15384 14977 15403 15011
rect 15403 14977 15436 15011
rect 15384 14968 15436 14977
rect 14740 14900 14792 14952
rect 15476 14900 15528 14952
rect 17960 14968 18012 15020
rect 18052 14968 18104 15020
rect 20260 15036 20312 15088
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 24676 15036 24728 15088
rect 21640 14968 21692 15020
rect 22376 14968 22428 15020
rect 24492 14968 24544 15020
rect 18696 14900 18748 14952
rect 18512 14832 18564 14884
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 19616 14943 19668 14952
rect 19616 14909 19625 14943
rect 19625 14909 19659 14943
rect 19659 14909 19668 14943
rect 19616 14900 19668 14909
rect 19800 14900 19852 14952
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 23388 14900 23440 14909
rect 19892 14832 19944 14884
rect 22008 14832 22060 14884
rect 22100 14832 22152 14884
rect 22376 14832 22428 14884
rect 24584 14832 24636 14884
rect 18420 14764 18472 14816
rect 20720 14764 20772 14816
rect 21916 14807 21968 14816
rect 21916 14773 21925 14807
rect 21925 14773 21959 14807
rect 21959 14773 21968 14807
rect 21916 14764 21968 14773
rect 25320 14764 25372 14816
rect 4043 14662 4095 14714
rect 4107 14662 4159 14714
rect 4171 14662 4223 14714
rect 4235 14662 4287 14714
rect 4299 14662 4351 14714
rect 10230 14662 10282 14714
rect 10294 14662 10346 14714
rect 10358 14662 10410 14714
rect 10422 14662 10474 14714
rect 10486 14662 10538 14714
rect 16417 14662 16469 14714
rect 16481 14662 16533 14714
rect 16545 14662 16597 14714
rect 16609 14662 16661 14714
rect 16673 14662 16725 14714
rect 22604 14662 22656 14714
rect 22668 14662 22720 14714
rect 22732 14662 22784 14714
rect 22796 14662 22848 14714
rect 22860 14662 22912 14714
rect 1860 14560 1912 14612
rect 2412 14560 2464 14612
rect 2964 14560 3016 14612
rect 940 14356 992 14408
rect 2872 14535 2924 14544
rect 2872 14501 2881 14535
rect 2881 14501 2915 14535
rect 2915 14501 2924 14535
rect 2872 14492 2924 14501
rect 5356 14535 5408 14544
rect 5356 14501 5365 14535
rect 5365 14501 5399 14535
rect 5399 14501 5408 14535
rect 5356 14492 5408 14501
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 3056 14424 3108 14476
rect 11888 14560 11940 14612
rect 14280 14560 14332 14612
rect 10048 14492 10100 14544
rect 6368 14424 6420 14476
rect 3884 14356 3936 14408
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 8208 14424 8260 14476
rect 15476 14424 15528 14476
rect 16672 14424 16724 14476
rect 4528 14288 4580 14340
rect 5080 14288 5132 14340
rect 3240 14220 3292 14272
rect 6000 14220 6052 14272
rect 6368 14288 6420 14340
rect 7840 14288 7892 14340
rect 8116 14288 8168 14340
rect 10508 14356 10560 14408
rect 14096 14356 14148 14408
rect 18052 14560 18104 14612
rect 19984 14560 20036 14612
rect 21916 14560 21968 14612
rect 18512 14535 18564 14544
rect 18512 14501 18521 14535
rect 18521 14501 18555 14535
rect 18555 14501 18564 14535
rect 18512 14492 18564 14501
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 19708 14356 19760 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 23388 14560 23440 14612
rect 23756 14560 23808 14612
rect 24492 14560 24544 14612
rect 25320 14560 25372 14612
rect 24584 14492 24636 14544
rect 24768 14492 24820 14544
rect 25964 14492 26016 14544
rect 10324 14288 10376 14340
rect 10784 14288 10836 14340
rect 11520 14288 11572 14340
rect 13636 14288 13688 14340
rect 15568 14288 15620 14340
rect 18420 14288 18472 14340
rect 21364 14288 21416 14340
rect 24860 14356 24912 14408
rect 24952 14356 25004 14408
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 8576 14220 8628 14272
rect 11612 14220 11664 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 15200 14220 15252 14272
rect 20536 14220 20588 14272
rect 24676 14288 24728 14340
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 4703 14118 4755 14170
rect 4767 14118 4819 14170
rect 4831 14118 4883 14170
rect 4895 14118 4947 14170
rect 4959 14118 5011 14170
rect 10890 14118 10942 14170
rect 10954 14118 11006 14170
rect 11018 14118 11070 14170
rect 11082 14118 11134 14170
rect 11146 14118 11198 14170
rect 17077 14118 17129 14170
rect 17141 14118 17193 14170
rect 17205 14118 17257 14170
rect 17269 14118 17321 14170
rect 17333 14118 17385 14170
rect 23264 14118 23316 14170
rect 23328 14118 23380 14170
rect 23392 14118 23444 14170
rect 23456 14118 23508 14170
rect 23520 14118 23572 14170
rect 3056 14016 3108 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 3240 14016 3292 14068
rect 4620 14016 4672 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 4436 13880 4488 13932
rect 5540 13948 5592 14000
rect 7104 14016 7156 14068
rect 6000 13880 6052 13932
rect 7380 13948 7432 14000
rect 10048 13948 10100 14000
rect 10324 14016 10376 14068
rect 10508 13948 10560 14000
rect 10784 13880 10836 13932
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 11796 13948 11848 14000
rect 12348 14016 12400 14068
rect 12532 14016 12584 14068
rect 12992 14016 13044 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 16304 14016 16356 14068
rect 21548 14016 21600 14068
rect 11612 13880 11664 13932
rect 3792 13855 3844 13864
rect 3792 13821 3801 13855
rect 3801 13821 3835 13855
rect 3835 13821 3844 13855
rect 3792 13812 3844 13821
rect 5080 13812 5132 13864
rect 5356 13812 5408 13864
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 9772 13812 9824 13864
rect 11244 13812 11296 13864
rect 11704 13812 11756 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 20996 13948 21048 14000
rect 24032 13991 24084 14000
rect 24032 13957 24041 13991
rect 24041 13957 24075 13991
rect 24075 13957 24084 13991
rect 24032 13948 24084 13957
rect 24492 13948 24544 14000
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 15292 13880 15344 13932
rect 14832 13812 14884 13864
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 16672 13880 16724 13932
rect 17960 13880 18012 13932
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 25504 13855 25556 13864
rect 25504 13821 25513 13855
rect 25513 13821 25547 13855
rect 25547 13821 25556 13855
rect 25504 13812 25556 13821
rect 6184 13744 6236 13796
rect 6552 13744 6604 13796
rect 8116 13744 8168 13796
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 5356 13719 5408 13728
rect 5356 13685 5365 13719
rect 5365 13685 5399 13719
rect 5399 13685 5408 13719
rect 5356 13676 5408 13685
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 8300 13676 8352 13728
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 10692 13787 10744 13796
rect 10692 13753 10701 13787
rect 10701 13753 10735 13787
rect 10735 13753 10744 13787
rect 10692 13744 10744 13753
rect 11612 13744 11664 13796
rect 12256 13744 12308 13796
rect 12164 13676 12216 13728
rect 12348 13719 12400 13728
rect 12348 13685 12357 13719
rect 12357 13685 12391 13719
rect 12391 13685 12400 13719
rect 12348 13676 12400 13685
rect 14280 13719 14332 13728
rect 14280 13685 14289 13719
rect 14289 13685 14323 13719
rect 14323 13685 14332 13719
rect 14280 13676 14332 13685
rect 14924 13744 14976 13796
rect 16856 13744 16908 13796
rect 17776 13744 17828 13796
rect 16764 13676 16816 13728
rect 17408 13676 17460 13728
rect 17868 13676 17920 13728
rect 4043 13574 4095 13626
rect 4107 13574 4159 13626
rect 4171 13574 4223 13626
rect 4235 13574 4287 13626
rect 4299 13574 4351 13626
rect 10230 13574 10282 13626
rect 10294 13574 10346 13626
rect 10358 13574 10410 13626
rect 10422 13574 10474 13626
rect 10486 13574 10538 13626
rect 16417 13574 16469 13626
rect 16481 13574 16533 13626
rect 16545 13574 16597 13626
rect 16609 13574 16661 13626
rect 16673 13574 16725 13626
rect 22604 13574 22656 13626
rect 22668 13574 22720 13626
rect 22732 13574 22784 13626
rect 22796 13574 22848 13626
rect 22860 13574 22912 13626
rect 7380 13472 7432 13524
rect 6184 13404 6236 13456
rect 7196 13447 7248 13456
rect 7196 13413 7205 13447
rect 7205 13413 7239 13447
rect 7239 13413 7248 13447
rect 7196 13404 7248 13413
rect 3792 13336 3844 13388
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 5080 13336 5132 13388
rect 5908 13336 5960 13388
rect 7012 13336 7064 13388
rect 3056 13200 3108 13252
rect 940 13132 992 13184
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 4528 13268 4580 13320
rect 5356 13268 5408 13320
rect 7196 13200 7248 13252
rect 8300 13404 8352 13456
rect 8760 13472 8812 13524
rect 10600 13472 10652 13524
rect 12532 13472 12584 13524
rect 12716 13472 12768 13524
rect 16672 13472 16724 13524
rect 16764 13472 16816 13524
rect 17684 13472 17736 13524
rect 18604 13472 18656 13524
rect 19984 13472 20036 13524
rect 20996 13515 21048 13524
rect 20996 13481 21005 13515
rect 21005 13481 21039 13515
rect 21039 13481 21048 13515
rect 20996 13472 21048 13481
rect 21364 13515 21416 13524
rect 21364 13481 21373 13515
rect 21373 13481 21407 13515
rect 21407 13481 21416 13515
rect 21364 13472 21416 13481
rect 24492 13515 24544 13524
rect 24492 13481 24501 13515
rect 24501 13481 24535 13515
rect 24535 13481 24544 13515
rect 24492 13472 24544 13481
rect 24860 13472 24912 13524
rect 8116 13379 8168 13388
rect 8116 13345 8125 13379
rect 8125 13345 8159 13379
rect 8159 13345 8168 13379
rect 8116 13336 8168 13345
rect 8392 13268 8444 13320
rect 4528 13132 4580 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 5080 13132 5132 13184
rect 5172 13132 5224 13184
rect 5356 13132 5408 13184
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 8116 13132 8168 13184
rect 9772 13336 9824 13388
rect 10048 13336 10100 13388
rect 12440 13336 12492 13388
rect 13636 13336 13688 13388
rect 17868 13336 17920 13388
rect 10784 13268 10836 13320
rect 10692 13200 10744 13252
rect 13452 13268 13504 13320
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 18052 13268 18104 13320
rect 12256 13200 12308 13252
rect 14280 13200 14332 13252
rect 15384 13200 15436 13252
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 12440 13132 12492 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 17408 13200 17460 13252
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 20260 13336 20312 13388
rect 20628 13336 20680 13388
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 18880 13200 18932 13252
rect 20536 13243 20588 13252
rect 20536 13209 20545 13243
rect 20545 13209 20579 13243
rect 20579 13209 20588 13243
rect 20536 13200 20588 13209
rect 25596 13268 25648 13320
rect 25688 13268 25740 13320
rect 18420 13175 18472 13184
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 18512 13132 18564 13184
rect 19340 13132 19392 13184
rect 21916 13132 21968 13184
rect 23664 13132 23716 13184
rect 25412 13175 25464 13184
rect 25412 13141 25421 13175
rect 25421 13141 25455 13175
rect 25455 13141 25464 13175
rect 25412 13132 25464 13141
rect 4703 13030 4755 13082
rect 4767 13030 4819 13082
rect 4831 13030 4883 13082
rect 4895 13030 4947 13082
rect 4959 13030 5011 13082
rect 10890 13030 10942 13082
rect 10954 13030 11006 13082
rect 11018 13030 11070 13082
rect 11082 13030 11134 13082
rect 11146 13030 11198 13082
rect 17077 13030 17129 13082
rect 17141 13030 17193 13082
rect 17205 13030 17257 13082
rect 17269 13030 17321 13082
rect 17333 13030 17385 13082
rect 23264 13030 23316 13082
rect 23328 13030 23380 13082
rect 23392 13030 23444 13082
rect 23456 13030 23508 13082
rect 23520 13030 23572 13082
rect 2872 12928 2924 12980
rect 4436 12928 4488 12980
rect 4712 12928 4764 12980
rect 6920 12928 6972 12980
rect 7564 12928 7616 12980
rect 8576 12928 8628 12980
rect 8668 12928 8720 12980
rect 10968 12928 11020 12980
rect 13268 12971 13320 12980
rect 4620 12860 4672 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 7656 12860 7708 12912
rect 8300 12860 8352 12912
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 13636 12928 13688 12980
rect 11244 12860 11296 12912
rect 14832 12860 14884 12912
rect 16120 12928 16172 12980
rect 16304 12928 16356 12980
rect 17960 12971 18012 12980
rect 17960 12937 17969 12971
rect 17969 12937 18003 12971
rect 18003 12937 18012 12971
rect 17960 12928 18012 12937
rect 21180 12928 21232 12980
rect 21548 12928 21600 12980
rect 15200 12903 15252 12912
rect 15200 12869 15209 12903
rect 15209 12869 15243 12903
rect 15243 12869 15252 12903
rect 15200 12860 15252 12869
rect 15292 12860 15344 12912
rect 16028 12860 16080 12912
rect 16580 12860 16632 12912
rect 18604 12860 18656 12912
rect 19340 12860 19392 12912
rect 20444 12860 20496 12912
rect 23112 12928 23164 12980
rect 23756 12928 23808 12980
rect 24400 12971 24452 12980
rect 24400 12937 24409 12971
rect 24409 12937 24443 12971
rect 24443 12937 24452 12971
rect 24400 12928 24452 12937
rect 24676 12928 24728 12980
rect 8116 12792 8168 12844
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 9772 12792 9824 12844
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 2136 12656 2188 12708
rect 2872 12588 2924 12640
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 5080 12724 5132 12776
rect 9680 12724 9732 12776
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 7840 12631 7892 12640
rect 7840 12597 7849 12631
rect 7849 12597 7883 12631
rect 7883 12597 7892 12631
rect 7840 12588 7892 12597
rect 9496 12656 9548 12708
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 11428 12792 11480 12844
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 12716 12792 12768 12844
rect 12992 12792 13044 12844
rect 12072 12724 12124 12776
rect 12348 12724 12400 12776
rect 9404 12588 9456 12640
rect 9864 12588 9916 12640
rect 11888 12656 11940 12708
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 10968 12588 11020 12640
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 12440 12588 12492 12640
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 17408 12792 17460 12844
rect 17868 12792 17920 12844
rect 20076 12835 20128 12844
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 15200 12724 15252 12776
rect 15752 12724 15804 12776
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 18880 12724 18932 12776
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 20260 12792 20312 12844
rect 23664 12860 23716 12912
rect 24584 12903 24636 12912
rect 24584 12869 24593 12903
rect 24593 12869 24627 12903
rect 24627 12869 24636 12903
rect 24584 12860 24636 12869
rect 26056 12792 26108 12844
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 20352 12724 20404 12776
rect 22928 12767 22980 12776
rect 22928 12733 22937 12767
rect 22937 12733 22971 12767
rect 22971 12733 22980 12767
rect 22928 12724 22980 12733
rect 13268 12656 13320 12708
rect 14924 12656 14976 12708
rect 17592 12588 17644 12640
rect 18052 12656 18104 12708
rect 20812 12656 20864 12708
rect 24860 12699 24912 12708
rect 24860 12665 24869 12699
rect 24869 12665 24903 12699
rect 24903 12665 24912 12699
rect 24860 12656 24912 12665
rect 25044 12656 25096 12708
rect 4043 12486 4095 12538
rect 4107 12486 4159 12538
rect 4171 12486 4223 12538
rect 4235 12486 4287 12538
rect 4299 12486 4351 12538
rect 10230 12486 10282 12538
rect 10294 12486 10346 12538
rect 10358 12486 10410 12538
rect 10422 12486 10474 12538
rect 10486 12486 10538 12538
rect 16417 12486 16469 12538
rect 16481 12486 16533 12538
rect 16545 12486 16597 12538
rect 16609 12486 16661 12538
rect 16673 12486 16725 12538
rect 22604 12486 22656 12538
rect 22668 12486 22720 12538
rect 22732 12486 22784 12538
rect 22796 12486 22848 12538
rect 22860 12486 22912 12538
rect 3056 12384 3108 12436
rect 3240 12384 3292 12436
rect 4896 12384 4948 12436
rect 2780 12316 2832 12368
rect 3884 12291 3936 12300
rect 3884 12257 3893 12291
rect 3893 12257 3927 12291
rect 3927 12257 3936 12291
rect 3884 12248 3936 12257
rect 4712 12248 4764 12300
rect 11520 12384 11572 12436
rect 12164 12384 12216 12436
rect 13636 12384 13688 12436
rect 15384 12384 15436 12436
rect 18328 12384 18380 12436
rect 19432 12384 19484 12436
rect 20352 12384 20404 12436
rect 23940 12384 23992 12436
rect 10876 12316 10928 12368
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 5540 12180 5592 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 8576 12248 8628 12300
rect 9404 12248 9456 12300
rect 10048 12248 10100 12300
rect 10692 12248 10744 12300
rect 13268 12359 13320 12368
rect 13268 12325 13277 12359
rect 13277 12325 13311 12359
rect 13311 12325 13320 12359
rect 13268 12316 13320 12325
rect 12992 12248 13044 12300
rect 2964 12112 3016 12164
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7840 12180 7892 12232
rect 9680 12180 9732 12232
rect 10784 12180 10836 12232
rect 12440 12180 12492 12232
rect 17408 12248 17460 12300
rect 17684 12248 17736 12300
rect 5816 12044 5868 12096
rect 11060 12112 11112 12164
rect 12164 12112 12216 12164
rect 13084 12112 13136 12164
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 11336 12044 11388 12096
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14464 12180 14516 12232
rect 18880 12359 18932 12368
rect 18880 12325 18889 12359
rect 18889 12325 18923 12359
rect 18923 12325 18932 12359
rect 18880 12316 18932 12325
rect 18604 12291 18656 12300
rect 18604 12257 18613 12291
rect 18613 12257 18647 12291
rect 18647 12257 18656 12291
rect 18604 12248 18656 12257
rect 18696 12248 18748 12300
rect 20536 12291 20588 12300
rect 20536 12257 20545 12291
rect 20545 12257 20579 12291
rect 20579 12257 20588 12291
rect 20536 12248 20588 12257
rect 21916 12316 21968 12368
rect 24032 12316 24084 12368
rect 24768 12316 24820 12368
rect 23848 12248 23900 12300
rect 24584 12248 24636 12300
rect 20444 12223 20496 12232
rect 20444 12189 20453 12223
rect 20453 12189 20487 12223
rect 20487 12189 20496 12223
rect 20444 12180 20496 12189
rect 23664 12180 23716 12232
rect 17684 12044 17736 12096
rect 17868 12044 17920 12096
rect 21456 12112 21508 12164
rect 22100 12112 22152 12164
rect 25964 12112 26016 12164
rect 4703 11942 4755 11994
rect 4767 11942 4819 11994
rect 4831 11942 4883 11994
rect 4895 11942 4947 11994
rect 4959 11942 5011 11994
rect 10890 11942 10942 11994
rect 10954 11942 11006 11994
rect 11018 11942 11070 11994
rect 11082 11942 11134 11994
rect 11146 11942 11198 11994
rect 17077 11942 17129 11994
rect 17141 11942 17193 11994
rect 17205 11942 17257 11994
rect 17269 11942 17321 11994
rect 17333 11942 17385 11994
rect 23264 11942 23316 11994
rect 23328 11942 23380 11994
rect 23392 11942 23444 11994
rect 23456 11942 23508 11994
rect 23520 11942 23572 11994
rect 2412 11883 2464 11892
rect 2412 11849 2421 11883
rect 2421 11849 2455 11883
rect 2455 11849 2464 11883
rect 2412 11840 2464 11849
rect 4528 11883 4580 11892
rect 4528 11849 4537 11883
rect 4537 11849 4571 11883
rect 4571 11849 4580 11883
rect 4528 11840 4580 11849
rect 3056 11815 3108 11824
rect 3056 11781 3065 11815
rect 3065 11781 3099 11815
rect 3099 11781 3108 11815
rect 3056 11772 3108 11781
rect 5080 11840 5132 11892
rect 6184 11840 6236 11892
rect 7564 11840 7616 11892
rect 8852 11840 8904 11892
rect 9588 11840 9640 11892
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 11520 11840 11572 11892
rect 11704 11840 11756 11892
rect 940 11704 992 11756
rect 1860 11636 1912 11688
rect 2780 11679 2832 11688
rect 1400 11568 1452 11620
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 5908 11704 5960 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 6828 11704 6880 11756
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 5080 11568 5132 11620
rect 7748 11704 7800 11756
rect 8208 11704 8260 11756
rect 20444 11840 20496 11892
rect 21456 11883 21508 11892
rect 21456 11849 21465 11883
rect 21465 11849 21499 11883
rect 21499 11849 21508 11883
rect 21456 11840 21508 11849
rect 9680 11772 9732 11824
rect 8300 11636 8352 11688
rect 6276 11568 6328 11620
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 11888 11704 11940 11756
rect 12072 11704 12124 11756
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10692 11500 10744 11552
rect 18328 11772 18380 11824
rect 20352 11772 20404 11824
rect 22376 11840 22428 11892
rect 23756 11840 23808 11892
rect 25136 11840 25188 11892
rect 25320 11840 25372 11892
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 17592 11704 17644 11756
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24768 11704 24820 11713
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 11612 11568 11664 11620
rect 11520 11500 11572 11552
rect 12164 11568 12216 11620
rect 18512 11568 18564 11620
rect 18788 11568 18840 11620
rect 20812 11568 20864 11620
rect 15844 11500 15896 11552
rect 17960 11500 18012 11552
rect 21364 11500 21416 11552
rect 23756 11636 23808 11688
rect 24400 11543 24452 11552
rect 24400 11509 24409 11543
rect 24409 11509 24443 11543
rect 24443 11509 24452 11543
rect 24400 11500 24452 11509
rect 4043 11398 4095 11450
rect 4107 11398 4159 11450
rect 4171 11398 4223 11450
rect 4235 11398 4287 11450
rect 4299 11398 4351 11450
rect 10230 11398 10282 11450
rect 10294 11398 10346 11450
rect 10358 11398 10410 11450
rect 10422 11398 10474 11450
rect 10486 11398 10538 11450
rect 16417 11398 16469 11450
rect 16481 11398 16533 11450
rect 16545 11398 16597 11450
rect 16609 11398 16661 11450
rect 16673 11398 16725 11450
rect 22604 11398 22656 11450
rect 22668 11398 22720 11450
rect 22732 11398 22784 11450
rect 22796 11398 22848 11450
rect 22860 11398 22912 11450
rect 3240 11160 3292 11212
rect 4528 11296 4580 11348
rect 6552 11296 6604 11348
rect 6828 11296 6880 11348
rect 7196 11339 7248 11348
rect 7196 11305 7205 11339
rect 7205 11305 7239 11339
rect 7239 11305 7248 11339
rect 9404 11339 9456 11348
rect 7196 11296 7248 11305
rect 8300 11271 8352 11280
rect 8300 11237 8309 11271
rect 8309 11237 8343 11271
rect 8343 11237 8352 11271
rect 8300 11228 8352 11237
rect 4528 11092 4580 11144
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 5724 11160 5776 11212
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 9404 11305 9434 11339
rect 9434 11305 9456 11339
rect 9404 11296 9456 11305
rect 10048 11296 10100 11348
rect 13728 11296 13780 11348
rect 14188 11296 14240 11348
rect 12624 11228 12676 11280
rect 13084 11228 13136 11280
rect 13912 11228 13964 11280
rect 14740 11296 14792 11348
rect 18880 11296 18932 11348
rect 22928 11296 22980 11348
rect 24400 11296 24452 11348
rect 24768 11296 24820 11348
rect 6552 11160 6604 11169
rect 2136 11024 2188 11076
rect 4160 11024 4212 11076
rect 6644 11092 6696 11144
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7288 11092 7340 11144
rect 7564 11024 7616 11076
rect 11336 11160 11388 11212
rect 11612 11160 11664 11212
rect 8668 11092 8720 11144
rect 8760 11092 8812 11144
rect 11060 11092 11112 11144
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 13360 11160 13412 11212
rect 15844 11160 15896 11212
rect 16212 11160 16264 11212
rect 14556 11092 14608 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 17960 11228 18012 11280
rect 17868 11203 17920 11212
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 5080 10956 5132 11008
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 16764 11024 16816 11076
rect 11060 10999 11112 11008
rect 11060 10965 11069 10999
rect 11069 10965 11103 10999
rect 11103 10965 11112 10999
rect 11060 10956 11112 10965
rect 11152 10956 11204 11008
rect 12440 10956 12492 11008
rect 14280 10956 14332 11008
rect 14740 10956 14792 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 16488 10999 16540 11008
rect 16488 10965 16497 10999
rect 16497 10965 16531 10999
rect 16531 10965 16540 10999
rect 16488 10956 16540 10965
rect 17316 11067 17368 11076
rect 17316 11033 17325 11067
rect 17325 11033 17359 11067
rect 17359 11033 17368 11067
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 20536 11160 20588 11212
rect 18696 11092 18748 11144
rect 18788 11092 18840 11144
rect 21180 11092 21232 11144
rect 24032 11271 24084 11280
rect 24032 11237 24041 11271
rect 24041 11237 24075 11271
rect 24075 11237 24084 11271
rect 24032 11228 24084 11237
rect 23664 11203 23716 11212
rect 23664 11169 23673 11203
rect 23673 11169 23707 11203
rect 23707 11169 23716 11203
rect 23664 11160 23716 11169
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 17316 11024 17368 11033
rect 21916 11024 21968 11076
rect 22100 11024 22152 11076
rect 25964 11024 26016 11076
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 21088 10999 21140 11008
rect 21088 10965 21097 10999
rect 21097 10965 21131 10999
rect 21131 10965 21140 10999
rect 21088 10956 21140 10965
rect 24400 10999 24452 11008
rect 24400 10965 24409 10999
rect 24409 10965 24443 10999
rect 24443 10965 24452 10999
rect 24400 10956 24452 10965
rect 24676 10999 24728 11008
rect 24676 10965 24685 10999
rect 24685 10965 24719 10999
rect 24719 10965 24728 10999
rect 24676 10956 24728 10965
rect 4703 10854 4755 10906
rect 4767 10854 4819 10906
rect 4831 10854 4883 10906
rect 4895 10854 4947 10906
rect 4959 10854 5011 10906
rect 10890 10854 10942 10906
rect 10954 10854 11006 10906
rect 11018 10854 11070 10906
rect 11082 10854 11134 10906
rect 11146 10854 11198 10906
rect 17077 10854 17129 10906
rect 17141 10854 17193 10906
rect 17205 10854 17257 10906
rect 17269 10854 17321 10906
rect 17333 10854 17385 10906
rect 23264 10854 23316 10906
rect 23328 10854 23380 10906
rect 23392 10854 23444 10906
rect 23456 10854 23508 10906
rect 23520 10854 23572 10906
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1860 10548 1912 10600
rect 4160 10616 4212 10668
rect 5540 10684 5592 10736
rect 5908 10684 5960 10736
rect 6644 10684 6696 10736
rect 7196 10684 7248 10736
rect 2320 10523 2372 10532
rect 2320 10489 2329 10523
rect 2329 10489 2363 10523
rect 2363 10489 2372 10523
rect 2320 10480 2372 10489
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 4804 10548 4856 10600
rect 5080 10616 5132 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 7104 10548 7156 10600
rect 8760 10752 8812 10804
rect 9680 10752 9732 10804
rect 10140 10752 10192 10804
rect 10784 10752 10836 10804
rect 11888 10752 11940 10804
rect 8484 10684 8536 10736
rect 12072 10684 12124 10736
rect 18052 10752 18104 10804
rect 18696 10752 18748 10804
rect 14004 10684 14056 10736
rect 9496 10616 9548 10668
rect 13544 10616 13596 10668
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 11980 10548 12032 10600
rect 13728 10616 13780 10668
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 16120 10616 16172 10668
rect 17224 10684 17276 10736
rect 18880 10752 18932 10804
rect 21088 10752 21140 10804
rect 24400 10752 24452 10804
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 23112 10616 23164 10668
rect 24676 10616 24728 10668
rect 25780 10616 25832 10668
rect 940 10412 992 10464
rect 2412 10412 2464 10464
rect 3516 10412 3568 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 6092 10480 6144 10532
rect 6552 10480 6604 10532
rect 6736 10480 6788 10532
rect 11612 10480 11664 10532
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 6828 10412 6880 10464
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 7748 10412 7800 10464
rect 12900 10412 12952 10464
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 14556 10412 14608 10464
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 17224 10548 17276 10600
rect 19800 10591 19852 10600
rect 19800 10557 19809 10591
rect 19809 10557 19843 10591
rect 19843 10557 19852 10591
rect 19800 10548 19852 10557
rect 23664 10548 23716 10600
rect 15844 10480 15896 10532
rect 16304 10480 16356 10532
rect 16488 10480 16540 10532
rect 16856 10480 16908 10532
rect 16212 10412 16264 10464
rect 21088 10412 21140 10464
rect 22284 10412 22336 10464
rect 23204 10455 23256 10464
rect 23204 10421 23213 10455
rect 23213 10421 23247 10455
rect 23247 10421 23256 10455
rect 23204 10412 23256 10421
rect 24032 10412 24084 10464
rect 24952 10412 25004 10464
rect 25412 10455 25464 10464
rect 25412 10421 25421 10455
rect 25421 10421 25455 10455
rect 25455 10421 25464 10455
rect 25412 10412 25464 10421
rect 4043 10310 4095 10362
rect 4107 10310 4159 10362
rect 4171 10310 4223 10362
rect 4235 10310 4287 10362
rect 4299 10310 4351 10362
rect 10230 10310 10282 10362
rect 10294 10310 10346 10362
rect 10358 10310 10410 10362
rect 10422 10310 10474 10362
rect 10486 10310 10538 10362
rect 16417 10310 16469 10362
rect 16481 10310 16533 10362
rect 16545 10310 16597 10362
rect 16609 10310 16661 10362
rect 16673 10310 16725 10362
rect 22604 10310 22656 10362
rect 22668 10310 22720 10362
rect 22732 10310 22784 10362
rect 22796 10310 22848 10362
rect 22860 10310 22912 10362
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 3516 10208 3568 10260
rect 4896 10208 4948 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7932 10208 7984 10260
rect 8484 10208 8536 10260
rect 11244 10208 11296 10260
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 6184 10140 6236 10192
rect 5908 10072 5960 10124
rect 11336 10140 11388 10192
rect 11980 10183 12032 10192
rect 11980 10149 11989 10183
rect 11989 10149 12023 10183
rect 12023 10149 12032 10183
rect 11980 10140 12032 10149
rect 11428 10072 11480 10124
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 13176 10208 13228 10260
rect 16028 10208 16080 10260
rect 13268 10140 13320 10192
rect 13084 10072 13136 10124
rect 2412 9936 2464 9988
rect 5356 10004 5408 10056
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3884 9868 3936 9920
rect 4804 9868 4856 9920
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 6920 9936 6972 9988
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 7932 10004 7984 10056
rect 8208 10004 8260 10056
rect 8392 10004 8444 10056
rect 9404 10004 9456 10056
rect 10140 10004 10192 10056
rect 11704 10004 11756 10056
rect 11888 10004 11940 10056
rect 12624 9979 12676 9988
rect 12624 9945 12633 9979
rect 12633 9945 12667 9979
rect 12667 9945 12676 9979
rect 12624 9936 12676 9945
rect 12716 9979 12768 9988
rect 12716 9945 12725 9979
rect 12725 9945 12759 9979
rect 12759 9945 12768 9979
rect 12716 9936 12768 9945
rect 13176 10004 13228 10056
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 14280 10004 14332 10056
rect 14924 10140 14976 10192
rect 14740 10115 14792 10124
rect 14740 10081 14749 10115
rect 14749 10081 14783 10115
rect 14783 10081 14792 10115
rect 14740 10072 14792 10081
rect 14648 10041 14700 10056
rect 15568 10140 15620 10192
rect 16856 10208 16908 10260
rect 17132 10208 17184 10260
rect 19892 10208 19944 10260
rect 22008 10208 22060 10260
rect 22744 10208 22796 10260
rect 23020 10208 23072 10260
rect 23204 10208 23256 10260
rect 16488 10072 16540 10124
rect 20628 10183 20680 10192
rect 20628 10149 20637 10183
rect 20637 10149 20671 10183
rect 20671 10149 20680 10183
rect 20628 10140 20680 10149
rect 21916 10140 21968 10192
rect 22376 10140 22428 10192
rect 14648 10007 14657 10041
rect 14657 10007 14691 10041
rect 14691 10007 14700 10041
rect 14648 10004 14700 10007
rect 15292 10004 15344 10056
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 16856 10004 16908 10056
rect 12900 9936 12952 9988
rect 13636 9936 13688 9988
rect 7932 9868 7984 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 10416 9911 10468 9920
rect 10416 9877 10425 9911
rect 10425 9877 10459 9911
rect 10459 9877 10468 9911
rect 10416 9868 10468 9877
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 12348 9868 12400 9920
rect 14096 9868 14148 9920
rect 15200 9936 15252 9988
rect 14832 9868 14884 9920
rect 15660 9868 15712 9920
rect 15844 9868 15896 9920
rect 16120 9868 16172 9920
rect 16488 9979 16540 9988
rect 16488 9945 16497 9979
rect 16497 9945 16531 9979
rect 16531 9945 16540 9979
rect 16488 9936 16540 9945
rect 16396 9868 16448 9920
rect 18420 10004 18472 10056
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 20352 10115 20404 10124
rect 20352 10081 20361 10115
rect 20361 10081 20395 10115
rect 20395 10081 20404 10115
rect 20352 10072 20404 10081
rect 21364 10072 21416 10124
rect 20720 10004 20772 10056
rect 25504 10208 25556 10260
rect 23756 10140 23808 10192
rect 24032 10140 24084 10192
rect 23664 10072 23716 10124
rect 24308 10004 24360 10056
rect 21180 9936 21232 9988
rect 21640 9936 21692 9988
rect 23020 9936 23072 9988
rect 17224 9868 17276 9920
rect 18788 9911 18840 9920
rect 18788 9877 18797 9911
rect 18797 9877 18831 9911
rect 18831 9877 18840 9911
rect 18788 9868 18840 9877
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 22468 9868 22520 9920
rect 23664 9911 23716 9920
rect 23664 9877 23673 9911
rect 23673 9877 23707 9911
rect 23707 9877 23716 9911
rect 23664 9868 23716 9877
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 4703 9766 4755 9818
rect 4767 9766 4819 9818
rect 4831 9766 4883 9818
rect 4895 9766 4947 9818
rect 4959 9766 5011 9818
rect 10890 9766 10942 9818
rect 10954 9766 11006 9818
rect 11018 9766 11070 9818
rect 11082 9766 11134 9818
rect 11146 9766 11198 9818
rect 17077 9766 17129 9818
rect 17141 9766 17193 9818
rect 17205 9766 17257 9818
rect 17269 9766 17321 9818
rect 17333 9766 17385 9818
rect 23264 9766 23316 9818
rect 23328 9766 23380 9818
rect 23392 9766 23444 9818
rect 23456 9766 23508 9818
rect 23520 9766 23572 9818
rect 25964 9732 26016 9784
rect 5448 9664 5500 9716
rect 6276 9664 6328 9716
rect 7840 9664 7892 9716
rect 3884 9528 3936 9580
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4712 9596 4764 9648
rect 7564 9596 7616 9648
rect 5540 9528 5592 9580
rect 5632 9528 5684 9580
rect 5724 9528 5776 9580
rect 6092 9528 6144 9580
rect 7012 9528 7064 9580
rect 7748 9528 7800 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 9312 9596 9364 9648
rect 10416 9596 10468 9648
rect 11704 9664 11756 9716
rect 11796 9664 11848 9716
rect 12164 9664 12216 9716
rect 12716 9664 12768 9716
rect 8392 9528 8444 9580
rect 8576 9528 8628 9580
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 3148 9460 3200 9512
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 940 9324 992 9376
rect 3148 9324 3200 9376
rect 11060 9460 11112 9512
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 12900 9596 12952 9648
rect 13176 9664 13228 9716
rect 13268 9639 13320 9648
rect 13268 9605 13293 9639
rect 13293 9605 13320 9639
rect 13268 9596 13320 9605
rect 12532 9571 12584 9580
rect 12532 9537 12550 9571
rect 12550 9537 12584 9571
rect 12532 9528 12584 9537
rect 10140 9392 10192 9444
rect 3700 9324 3752 9376
rect 4436 9324 4488 9376
rect 4620 9324 4672 9376
rect 7932 9324 7984 9376
rect 9772 9324 9824 9376
rect 10692 9324 10744 9376
rect 13084 9324 13136 9376
rect 17500 9664 17552 9716
rect 18052 9664 18104 9716
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13636 9528 13688 9580
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14832 9460 14884 9512
rect 15660 9528 15712 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 15292 9460 15344 9512
rect 16028 9528 16080 9580
rect 16488 9528 16540 9580
rect 19800 9596 19852 9648
rect 23112 9664 23164 9716
rect 23756 9664 23808 9716
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 20812 9528 20864 9580
rect 23664 9596 23716 9648
rect 16580 9460 16632 9512
rect 18788 9460 18840 9512
rect 22928 9503 22980 9512
rect 22928 9469 22937 9503
rect 22937 9469 22971 9503
rect 22971 9469 22980 9503
rect 22928 9460 22980 9469
rect 24860 9664 24912 9716
rect 24952 9707 25004 9716
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 24768 9460 24820 9512
rect 15476 9392 15528 9444
rect 15844 9392 15896 9444
rect 16672 9392 16724 9444
rect 17040 9392 17092 9444
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 15108 9324 15160 9376
rect 18328 9324 18380 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 24492 9367 24544 9376
rect 24492 9333 24501 9367
rect 24501 9333 24535 9367
rect 24535 9333 24544 9367
rect 24492 9324 24544 9333
rect 25320 9367 25372 9376
rect 25320 9333 25329 9367
rect 25329 9333 25363 9367
rect 25363 9333 25372 9367
rect 25320 9324 25372 9333
rect 4043 9222 4095 9274
rect 4107 9222 4159 9274
rect 4171 9222 4223 9274
rect 4235 9222 4287 9274
rect 4299 9222 4351 9274
rect 10230 9222 10282 9274
rect 10294 9222 10346 9274
rect 10358 9222 10410 9274
rect 10422 9222 10474 9274
rect 10486 9222 10538 9274
rect 16417 9222 16469 9274
rect 16481 9222 16533 9274
rect 16545 9222 16597 9274
rect 16609 9222 16661 9274
rect 16673 9222 16725 9274
rect 22604 9222 22656 9274
rect 22668 9222 22720 9274
rect 22732 9222 22784 9274
rect 22796 9222 22848 9274
rect 22860 9222 22912 9274
rect 3148 9120 3200 9172
rect 3332 9120 3384 9172
rect 4160 9052 4212 9104
rect 4712 9052 4764 9104
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 4436 8984 4488 9036
rect 4528 8984 4580 9036
rect 3424 8916 3476 8968
rect 3884 8916 3936 8968
rect 5540 9052 5592 9104
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 8300 9120 8352 9172
rect 8576 9052 8628 9104
rect 9772 9120 9824 9172
rect 9588 9052 9640 9104
rect 5356 8984 5408 9036
rect 6276 8984 6328 9036
rect 8668 8984 8720 9036
rect 11704 9052 11756 9104
rect 12348 9095 12400 9104
rect 12348 9061 12357 9095
rect 12357 9061 12391 9095
rect 12391 9061 12400 9095
rect 12348 9052 12400 9061
rect 11152 8984 11204 9036
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5816 8916 5868 8968
rect 9312 8916 9364 8968
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4436 8780 4488 8832
rect 8208 8848 8260 8900
rect 11244 8848 11296 8900
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 11980 8984 12032 9036
rect 13176 9120 13228 9172
rect 14188 9120 14240 9172
rect 14832 9120 14884 9172
rect 16028 9120 16080 9172
rect 20904 9120 20956 9172
rect 21180 9163 21232 9172
rect 21180 9129 21189 9163
rect 21189 9129 21223 9163
rect 21223 9129 21232 9163
rect 21180 9120 21232 9129
rect 22928 9120 22980 9172
rect 24492 9120 24544 9172
rect 12900 8984 12952 9036
rect 14004 9052 14056 9104
rect 15200 9052 15252 9104
rect 16856 9052 16908 9104
rect 17684 9052 17736 9104
rect 18696 8984 18748 9036
rect 19800 8984 19852 9036
rect 13544 8916 13596 8968
rect 14464 8916 14516 8968
rect 16028 8916 16080 8968
rect 16212 8959 16264 8968
rect 16212 8925 16221 8959
rect 16221 8925 16255 8959
rect 16255 8925 16264 8959
rect 16212 8916 16264 8925
rect 16672 8916 16724 8968
rect 17040 8916 17092 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 17960 8916 18012 8968
rect 19248 8916 19300 8968
rect 21272 8916 21324 8968
rect 24768 8984 24820 9036
rect 25228 8984 25280 9036
rect 5816 8780 5868 8832
rect 5908 8823 5960 8832
rect 5908 8789 5917 8823
rect 5917 8789 5951 8823
rect 5951 8789 5960 8823
rect 5908 8780 5960 8789
rect 9404 8780 9456 8832
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 15108 8848 15160 8900
rect 15660 8848 15712 8900
rect 14188 8780 14240 8832
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 21272 8823 21324 8832
rect 21272 8789 21281 8823
rect 21281 8789 21315 8823
rect 21315 8789 21324 8823
rect 21272 8780 21324 8789
rect 22008 8780 22060 8832
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 4703 8678 4755 8730
rect 4767 8678 4819 8730
rect 4831 8678 4883 8730
rect 4895 8678 4947 8730
rect 4959 8678 5011 8730
rect 10890 8678 10942 8730
rect 10954 8678 11006 8730
rect 11018 8678 11070 8730
rect 11082 8678 11134 8730
rect 11146 8678 11198 8730
rect 17077 8678 17129 8730
rect 17141 8678 17193 8730
rect 17205 8678 17257 8730
rect 17269 8678 17321 8730
rect 17333 8678 17385 8730
rect 23264 8678 23316 8730
rect 23328 8678 23380 8730
rect 23392 8678 23444 8730
rect 23456 8678 23508 8730
rect 23520 8678 23572 8730
rect 3792 8576 3844 8628
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 7840 8576 7892 8628
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 2044 8440 2096 8492
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3700 8483 3752 8492
rect 3700 8449 3718 8483
rect 3718 8449 3752 8483
rect 3700 8440 3752 8449
rect 3884 8440 3936 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4620 8440 4672 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 3424 8372 3476 8424
rect 4712 8372 4764 8424
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 9680 8551 9732 8560
rect 9680 8517 9689 8551
rect 9689 8517 9723 8551
rect 9723 8517 9732 8551
rect 9680 8508 9732 8517
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 8392 8440 8444 8492
rect 9588 8440 9640 8492
rect 10784 8508 10836 8560
rect 1676 8347 1728 8356
rect 1676 8313 1685 8347
rect 1685 8313 1719 8347
rect 1719 8313 1728 8347
rect 1676 8304 1728 8313
rect 2780 8304 2832 8356
rect 4344 8304 4396 8356
rect 12624 8576 12676 8628
rect 12900 8576 12952 8628
rect 11428 8440 11480 8492
rect 11980 8440 12032 8492
rect 12256 8508 12308 8560
rect 12716 8551 12768 8560
rect 12716 8517 12725 8551
rect 12725 8517 12759 8551
rect 12759 8517 12768 8551
rect 12716 8508 12768 8517
rect 14188 8619 14240 8628
rect 14188 8585 14197 8619
rect 14197 8585 14231 8619
rect 14231 8585 14240 8619
rect 14188 8576 14240 8585
rect 15660 8619 15712 8628
rect 15660 8585 15669 8619
rect 15669 8585 15703 8619
rect 15703 8585 15712 8619
rect 15660 8576 15712 8585
rect 16764 8576 16816 8628
rect 17684 8576 17736 8628
rect 18144 8576 18196 8628
rect 19892 8576 19944 8628
rect 20812 8619 20864 8628
rect 20812 8585 20821 8619
rect 20821 8585 20855 8619
rect 20855 8585 20864 8619
rect 20812 8576 20864 8585
rect 13820 8440 13872 8492
rect 12256 8372 12308 8424
rect 11704 8347 11756 8356
rect 11704 8313 11713 8347
rect 11713 8313 11747 8347
rect 11747 8313 11756 8347
rect 11704 8304 11756 8313
rect 18052 8508 18104 8560
rect 20352 8551 20404 8560
rect 20352 8517 20361 8551
rect 20361 8517 20395 8551
rect 20395 8517 20404 8551
rect 20352 8508 20404 8517
rect 25320 8508 25372 8560
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 17500 8415 17552 8424
rect 17500 8381 17509 8415
rect 17509 8381 17543 8415
rect 17543 8381 17552 8415
rect 17500 8372 17552 8381
rect 18696 8372 18748 8424
rect 20720 8372 20772 8424
rect 20628 8347 20680 8356
rect 20628 8313 20637 8347
rect 20637 8313 20671 8347
rect 20671 8313 20680 8347
rect 20628 8304 20680 8313
rect 1952 8279 2004 8288
rect 1952 8245 1961 8279
rect 1961 8245 1995 8279
rect 1995 8245 2004 8279
rect 1952 8236 2004 8245
rect 3516 8279 3568 8288
rect 3516 8245 3525 8279
rect 3525 8245 3559 8279
rect 3559 8245 3568 8279
rect 3516 8236 3568 8245
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 7840 8236 7892 8288
rect 12164 8236 12216 8288
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 18052 8236 18104 8288
rect 22008 8304 22060 8356
rect 25228 8304 25280 8356
rect 25872 8304 25924 8356
rect 22100 8236 22152 8288
rect 22192 8236 22244 8288
rect 23112 8236 23164 8288
rect 4043 8134 4095 8186
rect 4107 8134 4159 8186
rect 4171 8134 4223 8186
rect 4235 8134 4287 8186
rect 4299 8134 4351 8186
rect 10230 8134 10282 8186
rect 10294 8134 10346 8186
rect 10358 8134 10410 8186
rect 10422 8134 10474 8186
rect 10486 8134 10538 8186
rect 16417 8134 16469 8186
rect 16481 8134 16533 8186
rect 16545 8134 16597 8186
rect 16609 8134 16661 8186
rect 16673 8134 16725 8186
rect 22604 8134 22656 8186
rect 22668 8134 22720 8186
rect 22732 8134 22784 8186
rect 22796 8134 22848 8186
rect 22860 8134 22912 8186
rect 3792 8032 3844 8084
rect 7380 8032 7432 8084
rect 7656 8032 7708 8084
rect 8760 8032 8812 8084
rect 9772 8032 9824 8084
rect 13820 8032 13872 8084
rect 13912 8032 13964 8084
rect 16212 8032 16264 8084
rect 17960 8075 18012 8084
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 18420 8032 18472 8084
rect 4436 7964 4488 8016
rect 6092 7964 6144 8016
rect 3516 7896 3568 7948
rect 2780 7828 2832 7880
rect 4804 7896 4856 7948
rect 5816 7896 5868 7948
rect 6920 7896 6972 7948
rect 1952 7760 2004 7812
rect 4620 7828 4672 7880
rect 5908 7828 5960 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 3056 7692 3108 7744
rect 4712 7760 4764 7812
rect 6092 7760 6144 7812
rect 3608 7692 3660 7744
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 8208 7964 8260 8016
rect 8668 8007 8720 8016
rect 8668 7973 8677 8007
rect 8677 7973 8711 8007
rect 8711 7973 8720 8007
rect 8668 7964 8720 7973
rect 11244 7964 11296 8016
rect 12256 7964 12308 8016
rect 13360 7964 13412 8016
rect 7472 7896 7524 7948
rect 8300 7896 8352 7948
rect 7748 7828 7800 7880
rect 8484 7828 8536 7880
rect 8852 7828 8904 7880
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 11888 7760 11940 7812
rect 7104 7692 7156 7744
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 8208 7692 8260 7744
rect 8944 7692 8996 7744
rect 11612 7692 11664 7744
rect 14188 7692 14240 7744
rect 17500 7964 17552 8016
rect 17776 8007 17828 8016
rect 17776 7973 17785 8007
rect 17785 7973 17819 8007
rect 17819 7973 17828 8007
rect 17776 7964 17828 7973
rect 17224 7896 17276 7948
rect 16580 7828 16632 7880
rect 17868 7828 17920 7880
rect 22192 7964 22244 8016
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 21180 7896 21232 7948
rect 15016 7760 15068 7812
rect 15568 7760 15620 7812
rect 17776 7760 17828 7812
rect 20720 7828 20772 7880
rect 22100 7828 22152 7880
rect 18420 7760 18472 7812
rect 25964 7828 26016 7880
rect 17684 7692 17736 7744
rect 19248 7692 19300 7744
rect 22100 7692 22152 7744
rect 24952 7692 25004 7744
rect 25688 7692 25740 7744
rect 4703 7590 4755 7642
rect 4767 7590 4819 7642
rect 4831 7590 4883 7642
rect 4895 7590 4947 7642
rect 4959 7590 5011 7642
rect 10890 7590 10942 7642
rect 10954 7590 11006 7642
rect 11018 7590 11070 7642
rect 11082 7590 11134 7642
rect 11146 7590 11198 7642
rect 17077 7590 17129 7642
rect 17141 7590 17193 7642
rect 17205 7590 17257 7642
rect 17269 7590 17321 7642
rect 17333 7590 17385 7642
rect 23264 7590 23316 7642
rect 23328 7590 23380 7642
rect 23392 7590 23444 7642
rect 23456 7590 23508 7642
rect 23520 7590 23572 7642
rect 940 7488 992 7540
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2044 7420 2096 7472
rect 7104 7488 7156 7540
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 7012 7420 7064 7472
rect 2780 7352 2832 7404
rect 6092 7395 6144 7404
rect 6092 7361 6101 7395
rect 6101 7361 6135 7395
rect 6135 7361 6144 7395
rect 6092 7352 6144 7361
rect 8392 7488 8444 7540
rect 8576 7488 8628 7540
rect 8668 7488 8720 7540
rect 8944 7488 8996 7540
rect 7748 7420 7800 7472
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 5816 7284 5868 7336
rect 2412 7259 2464 7268
rect 2412 7225 2421 7259
rect 2421 7225 2455 7259
rect 2455 7225 2464 7259
rect 2412 7216 2464 7225
rect 4620 7148 4672 7200
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 7840 7259 7892 7268
rect 7840 7225 7849 7259
rect 7849 7225 7883 7259
rect 7883 7225 7892 7259
rect 7840 7216 7892 7225
rect 8300 7259 8352 7268
rect 8300 7225 8309 7259
rect 8309 7225 8343 7259
rect 8343 7225 8352 7259
rect 8300 7216 8352 7225
rect 6368 7148 6420 7200
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 7748 7148 7800 7200
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9036 7352 9088 7404
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 9312 7420 9364 7472
rect 9680 7463 9732 7472
rect 9680 7429 9705 7463
rect 9705 7429 9732 7463
rect 9680 7420 9732 7429
rect 12440 7420 12492 7472
rect 12624 7488 12676 7540
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 14096 7420 14148 7472
rect 16580 7488 16632 7540
rect 16948 7488 17000 7540
rect 17960 7488 18012 7540
rect 18512 7488 18564 7540
rect 20996 7488 21048 7540
rect 16212 7420 16264 7472
rect 15660 7352 15712 7404
rect 22192 7463 22244 7472
rect 22192 7429 22201 7463
rect 22201 7429 22235 7463
rect 22235 7429 22244 7463
rect 22192 7420 22244 7429
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 11980 7284 12032 7336
rect 12072 7284 12124 7336
rect 12256 7284 12308 7336
rect 15936 7284 15988 7336
rect 16304 7284 16356 7336
rect 18052 7352 18104 7404
rect 18144 7352 18196 7404
rect 18512 7395 18564 7404
rect 18512 7361 18521 7395
rect 18521 7361 18555 7395
rect 18555 7361 18564 7395
rect 18512 7352 18564 7361
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 19892 7352 19944 7404
rect 11888 7216 11940 7268
rect 13452 7216 13504 7268
rect 15108 7216 15160 7268
rect 15384 7259 15436 7268
rect 15384 7225 15393 7259
rect 15393 7225 15427 7259
rect 15427 7225 15436 7259
rect 15384 7216 15436 7225
rect 18328 7284 18380 7336
rect 8668 7148 8720 7200
rect 9128 7148 9180 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 11612 7148 11664 7200
rect 15016 7148 15068 7200
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 17408 7216 17460 7268
rect 23112 7420 23164 7472
rect 17684 7148 17736 7200
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 19340 7148 19392 7200
rect 21180 7191 21232 7200
rect 21180 7157 21189 7191
rect 21189 7157 21223 7191
rect 21223 7157 21232 7191
rect 21180 7148 21232 7157
rect 4043 7046 4095 7098
rect 4107 7046 4159 7098
rect 4171 7046 4223 7098
rect 4235 7046 4287 7098
rect 4299 7046 4351 7098
rect 10230 7046 10282 7098
rect 10294 7046 10346 7098
rect 10358 7046 10410 7098
rect 10422 7046 10474 7098
rect 10486 7046 10538 7098
rect 16417 7046 16469 7098
rect 16481 7046 16533 7098
rect 16545 7046 16597 7098
rect 16609 7046 16661 7098
rect 16673 7046 16725 7098
rect 22604 7046 22656 7098
rect 22668 7046 22720 7098
rect 22732 7046 22784 7098
rect 22796 7046 22848 7098
rect 22860 7046 22912 7098
rect 7840 6944 7892 6996
rect 2412 6808 2464 6860
rect 4712 6876 4764 6928
rect 6092 6876 6144 6928
rect 6828 6876 6880 6928
rect 8668 6944 8720 6996
rect 8852 6944 8904 6996
rect 9128 6944 9180 6996
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 3792 6740 3844 6792
rect 5356 6740 5408 6792
rect 6276 6808 6328 6860
rect 2044 6672 2096 6724
rect 8760 6808 8812 6860
rect 6920 6740 6972 6792
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7472 6672 7524 6724
rect 5356 6604 5408 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 7840 6604 7892 6656
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8484 6740 8536 6792
rect 9404 6919 9456 6928
rect 9404 6885 9413 6919
rect 9413 6885 9447 6919
rect 9447 6885 9456 6919
rect 9404 6876 9456 6885
rect 12440 6944 12492 6996
rect 14280 6944 14332 6996
rect 15016 6944 15068 6996
rect 18052 6944 18104 6996
rect 18512 6944 18564 6996
rect 18972 6944 19024 6996
rect 25964 6944 26016 6996
rect 10784 6876 10836 6928
rect 8300 6715 8352 6724
rect 8300 6681 8309 6715
rect 8309 6681 8343 6715
rect 8343 6681 8352 6715
rect 9128 6740 9180 6792
rect 9312 6740 9364 6792
rect 15384 6876 15436 6928
rect 17960 6919 18012 6928
rect 17960 6885 17969 6919
rect 17969 6885 18003 6919
rect 18003 6885 18012 6919
rect 17960 6876 18012 6885
rect 11336 6808 11388 6860
rect 12072 6808 12124 6860
rect 12256 6808 12308 6860
rect 19800 6808 19852 6860
rect 22376 6808 22428 6860
rect 8300 6672 8352 6681
rect 9036 6672 9088 6724
rect 9404 6672 9456 6724
rect 9772 6740 9824 6792
rect 11244 6740 11296 6792
rect 16212 6740 16264 6792
rect 16948 6740 17000 6792
rect 17776 6740 17828 6792
rect 18052 6740 18104 6792
rect 18972 6740 19024 6792
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 9680 6604 9732 6656
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 12348 6672 12400 6724
rect 15660 6672 15712 6724
rect 16304 6672 16356 6724
rect 19248 6672 19300 6724
rect 11888 6604 11940 6656
rect 16120 6604 16172 6656
rect 20076 6604 20128 6656
rect 20812 6715 20864 6724
rect 20812 6681 20821 6715
rect 20821 6681 20855 6715
rect 20855 6681 20864 6715
rect 20812 6672 20864 6681
rect 21456 6672 21508 6724
rect 20720 6604 20772 6656
rect 21732 6604 21784 6656
rect 4703 6502 4755 6554
rect 4767 6502 4819 6554
rect 4831 6502 4883 6554
rect 4895 6502 4947 6554
rect 4959 6502 5011 6554
rect 10890 6502 10942 6554
rect 10954 6502 11006 6554
rect 11018 6502 11070 6554
rect 11082 6502 11134 6554
rect 11146 6502 11198 6554
rect 17077 6502 17129 6554
rect 17141 6502 17193 6554
rect 17205 6502 17257 6554
rect 17269 6502 17321 6554
rect 17333 6502 17385 6554
rect 23264 6502 23316 6554
rect 23328 6502 23380 6554
rect 23392 6502 23444 6554
rect 23456 6502 23508 6554
rect 23520 6502 23572 6554
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4712 6307 4764 6316
rect 4712 6273 4721 6307
rect 4721 6273 4755 6307
rect 4755 6273 4764 6307
rect 4712 6264 4764 6273
rect 5356 6264 5408 6316
rect 2688 6196 2740 6248
rect 7012 6400 7064 6452
rect 7196 6400 7248 6452
rect 7748 6400 7800 6452
rect 8300 6400 8352 6452
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6184 6264 6236 6316
rect 7012 6264 7064 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 4620 6060 4672 6112
rect 5080 6060 5132 6112
rect 5264 6060 5316 6112
rect 6736 6060 6788 6112
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 7656 6060 7708 6112
rect 8392 6332 8444 6384
rect 8760 6400 8812 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 9220 6400 9272 6452
rect 9680 6400 9732 6452
rect 11704 6400 11756 6452
rect 11888 6400 11940 6452
rect 12348 6443 12400 6452
rect 12348 6409 12357 6443
rect 12357 6409 12391 6443
rect 12391 6409 12400 6443
rect 12348 6400 12400 6409
rect 14832 6443 14884 6452
rect 14832 6409 14841 6443
rect 14841 6409 14875 6443
rect 14875 6409 14884 6443
rect 14832 6400 14884 6409
rect 15660 6400 15712 6452
rect 15844 6400 15896 6452
rect 16304 6400 16356 6452
rect 16396 6400 16448 6452
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 11612 6332 11664 6384
rect 14096 6332 14148 6384
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 10692 6264 10744 6316
rect 9680 6128 9732 6180
rect 12072 6171 12124 6180
rect 12072 6137 12081 6171
rect 12081 6137 12115 6171
rect 12115 6137 12124 6171
rect 12072 6128 12124 6137
rect 12164 6128 12216 6180
rect 13912 6128 13964 6180
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 18052 6332 18104 6384
rect 18328 6375 18380 6384
rect 18328 6341 18337 6375
rect 18337 6341 18371 6375
rect 18371 6341 18380 6375
rect 18328 6332 18380 6341
rect 19340 6332 19392 6384
rect 19800 6443 19852 6452
rect 19800 6409 19809 6443
rect 19809 6409 19843 6443
rect 19843 6409 19852 6443
rect 19800 6400 19852 6409
rect 20812 6400 20864 6452
rect 21456 6443 21508 6452
rect 21456 6409 21465 6443
rect 21465 6409 21499 6443
rect 21499 6409 21508 6443
rect 21456 6400 21508 6409
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 14372 6128 14424 6180
rect 10232 6060 10284 6112
rect 11428 6060 11480 6112
rect 13636 6060 13688 6112
rect 14832 6060 14884 6112
rect 15016 6128 15068 6180
rect 15568 6128 15620 6180
rect 15752 6196 15804 6248
rect 16304 6307 16356 6316
rect 16304 6273 16318 6307
rect 16318 6273 16352 6307
rect 16352 6273 16356 6307
rect 16304 6264 16356 6273
rect 20352 6264 20404 6316
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 17316 6196 17368 6248
rect 17684 6128 17736 6180
rect 17960 6128 18012 6180
rect 16396 6060 16448 6112
rect 17132 6103 17184 6112
rect 17132 6069 17141 6103
rect 17141 6069 17175 6103
rect 17175 6069 17184 6103
rect 17132 6060 17184 6069
rect 18420 6196 18472 6248
rect 20444 6128 20496 6180
rect 21732 6264 21784 6316
rect 25504 6264 25556 6316
rect 24124 6128 24176 6180
rect 25412 6171 25464 6180
rect 25412 6137 25421 6171
rect 25421 6137 25455 6171
rect 25455 6137 25464 6171
rect 25412 6128 25464 6137
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 22376 6060 22428 6112
rect 22836 6060 22888 6112
rect 4043 5958 4095 6010
rect 4107 5958 4159 6010
rect 4171 5958 4223 6010
rect 4235 5958 4287 6010
rect 4299 5958 4351 6010
rect 10230 5958 10282 6010
rect 10294 5958 10346 6010
rect 10358 5958 10410 6010
rect 10422 5958 10474 6010
rect 10486 5958 10538 6010
rect 16417 5958 16469 6010
rect 16481 5958 16533 6010
rect 16545 5958 16597 6010
rect 16609 5958 16661 6010
rect 16673 5958 16725 6010
rect 22604 5958 22656 6010
rect 22668 5958 22720 6010
rect 22732 5958 22784 6010
rect 22796 5958 22848 6010
rect 22860 5958 22912 6010
rect 7380 5856 7432 5908
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 7564 5856 7616 5908
rect 6736 5788 6788 5840
rect 5264 5720 5316 5772
rect 7012 5763 7064 5772
rect 7012 5729 7021 5763
rect 7021 5729 7055 5763
rect 7055 5729 7064 5763
rect 7012 5720 7064 5729
rect 7656 5788 7708 5840
rect 8760 5856 8812 5908
rect 11336 5856 11388 5908
rect 13912 5856 13964 5908
rect 9404 5788 9456 5840
rect 4436 5652 4488 5704
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 5448 5584 5500 5636
rect 7380 5584 7432 5636
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 15200 5856 15252 5908
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 15660 5788 15712 5840
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 15752 5763 15804 5772
rect 13636 5584 13688 5636
rect 14372 5652 14424 5704
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 16948 5856 17000 5908
rect 17224 5856 17276 5908
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 14280 5584 14332 5636
rect 8944 5516 8996 5568
rect 12440 5516 12492 5568
rect 15292 5584 15344 5636
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 17132 5788 17184 5840
rect 19800 5856 19852 5908
rect 21732 5856 21784 5908
rect 20444 5788 20496 5840
rect 20720 5788 20772 5840
rect 16212 5652 16264 5704
rect 17132 5652 17184 5704
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 18052 5652 18104 5704
rect 20352 5763 20404 5772
rect 20352 5729 20361 5763
rect 20361 5729 20395 5763
rect 20395 5729 20404 5763
rect 20352 5720 20404 5729
rect 21180 5763 21232 5772
rect 21180 5729 21189 5763
rect 21189 5729 21223 5763
rect 21223 5729 21232 5763
rect 21180 5720 21232 5729
rect 19524 5652 19576 5704
rect 20536 5652 20588 5704
rect 15660 5516 15712 5568
rect 16488 5516 16540 5568
rect 20076 5584 20128 5636
rect 21824 5584 21876 5636
rect 23112 5516 23164 5568
rect 4703 5414 4755 5466
rect 4767 5414 4819 5466
rect 4831 5414 4883 5466
rect 4895 5414 4947 5466
rect 4959 5414 5011 5466
rect 10890 5414 10942 5466
rect 10954 5414 11006 5466
rect 11018 5414 11070 5466
rect 11082 5414 11134 5466
rect 11146 5414 11198 5466
rect 17077 5414 17129 5466
rect 17141 5414 17193 5466
rect 17205 5414 17257 5466
rect 17269 5414 17321 5466
rect 17333 5414 17385 5466
rect 23264 5414 23316 5466
rect 23328 5414 23380 5466
rect 23392 5414 23444 5466
rect 23456 5414 23508 5466
rect 23520 5414 23572 5466
rect 4436 5312 4488 5364
rect 5080 5312 5132 5364
rect 940 5176 992 5228
rect 6828 5312 6880 5364
rect 7656 5176 7708 5228
rect 7932 5312 7984 5364
rect 8392 5312 8444 5364
rect 9496 5244 9548 5296
rect 12440 5244 12492 5296
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 14004 5312 14056 5364
rect 14464 5176 14516 5228
rect 4620 5108 4672 5160
rect 11244 5108 11296 5160
rect 14832 5176 14884 5228
rect 15292 5176 15344 5228
rect 15476 5182 15528 5234
rect 16764 5312 16816 5364
rect 16948 5312 17000 5364
rect 17868 5312 17920 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 20812 5312 20864 5364
rect 17408 5244 17460 5296
rect 18236 5287 18288 5296
rect 18236 5253 18245 5287
rect 18245 5253 18279 5287
rect 18279 5253 18288 5287
rect 18236 5244 18288 5253
rect 20352 5244 20404 5296
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 15568 5108 15620 5160
rect 16028 5176 16080 5228
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 18788 5176 18840 5228
rect 20352 5108 20404 5160
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 22100 5176 22152 5228
rect 23020 5176 23072 5228
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 21732 5108 21784 5160
rect 20444 5083 20496 5092
rect 20444 5049 20453 5083
rect 20453 5049 20487 5083
rect 20487 5049 20496 5083
rect 20444 5040 20496 5049
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 8024 4972 8076 5024
rect 9036 4972 9088 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 14096 4972 14148 5024
rect 14924 5015 14976 5024
rect 14924 4981 14933 5015
rect 14933 4981 14967 5015
rect 14967 4981 14976 5015
rect 14924 4972 14976 4981
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 16028 4972 16080 5024
rect 16120 4972 16172 5024
rect 16304 4972 16356 5024
rect 20628 5015 20680 5024
rect 20628 4981 20637 5015
rect 20637 4981 20671 5015
rect 20671 4981 20680 5015
rect 20628 4972 20680 4981
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 4043 4870 4095 4922
rect 4107 4870 4159 4922
rect 4171 4870 4223 4922
rect 4235 4870 4287 4922
rect 4299 4870 4351 4922
rect 10230 4870 10282 4922
rect 10294 4870 10346 4922
rect 10358 4870 10410 4922
rect 10422 4870 10474 4922
rect 10486 4870 10538 4922
rect 16417 4870 16469 4922
rect 16481 4870 16533 4922
rect 16545 4870 16597 4922
rect 16609 4870 16661 4922
rect 16673 4870 16725 4922
rect 22604 4870 22656 4922
rect 22668 4870 22720 4922
rect 22732 4870 22784 4922
rect 22796 4870 22848 4922
rect 22860 4870 22912 4922
rect 940 4564 992 4616
rect 5724 4564 5776 4616
rect 7656 4768 7708 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8024 4564 8076 4616
rect 11336 4768 11388 4820
rect 13820 4768 13872 4820
rect 12164 4700 12216 4752
rect 12716 4700 12768 4752
rect 9772 4564 9824 4616
rect 10692 4632 10744 4684
rect 12256 4632 12308 4684
rect 12900 4632 12952 4684
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 14280 4700 14332 4752
rect 15752 4768 15804 4820
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 16304 4811 16356 4820
rect 16304 4777 16313 4811
rect 16313 4777 16347 4811
rect 16347 4777 16356 4811
rect 16304 4768 16356 4777
rect 19248 4768 19300 4820
rect 20628 4768 20680 4820
rect 14924 4700 14976 4752
rect 14648 4632 14700 4684
rect 11980 4564 12032 4616
rect 15752 4632 15804 4684
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 15568 4564 15620 4616
rect 15660 4564 15712 4616
rect 16396 4700 16448 4752
rect 16764 4564 16816 4616
rect 17868 4632 17920 4684
rect 23112 4564 23164 4616
rect 25228 4607 25280 4616
rect 25228 4573 25237 4607
rect 25237 4573 25271 4607
rect 25271 4573 25280 4607
rect 25228 4564 25280 4573
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 7564 4428 7616 4480
rect 15476 4496 15528 4548
rect 17960 4496 18012 4548
rect 10324 4428 10376 4480
rect 13912 4428 13964 4480
rect 15844 4428 15896 4480
rect 20904 4428 20956 4480
rect 22100 4428 22152 4480
rect 25412 4471 25464 4480
rect 25412 4437 25421 4471
rect 25421 4437 25455 4471
rect 25455 4437 25464 4471
rect 25412 4428 25464 4437
rect 4703 4326 4755 4378
rect 4767 4326 4819 4378
rect 4831 4326 4883 4378
rect 4895 4326 4947 4378
rect 4959 4326 5011 4378
rect 10890 4326 10942 4378
rect 10954 4326 11006 4378
rect 11018 4326 11070 4378
rect 11082 4326 11134 4378
rect 11146 4326 11198 4378
rect 17077 4326 17129 4378
rect 17141 4326 17193 4378
rect 17205 4326 17257 4378
rect 17269 4326 17321 4378
rect 17333 4326 17385 4378
rect 23264 4326 23316 4378
rect 23328 4326 23380 4378
rect 23392 4326 23444 4378
rect 23456 4326 23508 4378
rect 23520 4326 23572 4378
rect 5448 4224 5500 4276
rect 11980 4224 12032 4276
rect 14280 4224 14332 4276
rect 14740 4267 14792 4276
rect 14740 4233 14749 4267
rect 14749 4233 14783 4267
rect 14783 4233 14792 4267
rect 14740 4224 14792 4233
rect 14832 4224 14884 4276
rect 17960 4224 18012 4276
rect 22284 4224 22336 4276
rect 7932 4156 7984 4208
rect 9588 4156 9640 4208
rect 10324 4156 10376 4208
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 6000 4020 6052 4072
rect 7380 4088 7432 4140
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 7840 4088 7892 4140
rect 8024 4088 8076 4140
rect 11060 4131 11112 4140
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 8208 4020 8260 4072
rect 8300 4020 8352 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 7932 3952 7984 4004
rect 6000 3927 6052 3936
rect 6000 3893 6009 3927
rect 6009 3893 6043 3927
rect 6043 3893 6052 3927
rect 6000 3884 6052 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 8944 3952 8996 4004
rect 10784 3995 10836 4004
rect 10784 3961 10793 3995
rect 10793 3961 10827 3995
rect 10827 3961 10836 3995
rect 10784 3952 10836 3961
rect 12716 4020 12768 4072
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 20904 4156 20956 4208
rect 15292 4088 15344 4140
rect 15016 4020 15068 4072
rect 17684 4088 17736 4140
rect 19524 4088 19576 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 19708 4020 19760 4072
rect 12900 3995 12952 4004
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 13728 3995 13780 4004
rect 13728 3961 13737 3995
rect 13737 3961 13771 3995
rect 13771 3961 13780 3995
rect 13728 3952 13780 3961
rect 15660 3952 15712 4004
rect 17500 3952 17552 4004
rect 8392 3884 8444 3936
rect 9864 3884 9916 3936
rect 12624 3884 12676 3936
rect 14280 3884 14332 3936
rect 22284 3884 22336 3936
rect 23664 3884 23716 3936
rect 24952 3884 25004 3936
rect 4043 3782 4095 3834
rect 4107 3782 4159 3834
rect 4171 3782 4223 3834
rect 4235 3782 4287 3834
rect 4299 3782 4351 3834
rect 10230 3782 10282 3834
rect 10294 3782 10346 3834
rect 10358 3782 10410 3834
rect 10422 3782 10474 3834
rect 10486 3782 10538 3834
rect 16417 3782 16469 3834
rect 16481 3782 16533 3834
rect 16545 3782 16597 3834
rect 16609 3782 16661 3834
rect 16673 3782 16725 3834
rect 22604 3782 22656 3834
rect 22668 3782 22720 3834
rect 22732 3782 22784 3834
rect 22796 3782 22848 3834
rect 22860 3782 22912 3834
rect 5264 3680 5316 3732
rect 7012 3680 7064 3732
rect 7380 3680 7432 3732
rect 8208 3680 8260 3732
rect 11060 3680 11112 3732
rect 11428 3680 11480 3732
rect 7840 3655 7892 3664
rect 7840 3621 7849 3655
rect 7849 3621 7883 3655
rect 7883 3621 7892 3655
rect 7840 3612 7892 3621
rect 1032 3476 1084 3528
rect 8300 3544 8352 3596
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 7748 3476 7800 3528
rect 10692 3544 10744 3596
rect 11244 3544 11296 3596
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 4436 3408 4488 3460
rect 4528 3451 4580 3460
rect 4528 3417 4537 3451
rect 4537 3417 4571 3451
rect 4571 3417 4580 3451
rect 4528 3408 4580 3417
rect 4620 3408 4672 3460
rect 5816 3408 5868 3460
rect 7104 3408 7156 3460
rect 9128 3408 9180 3460
rect 9588 3408 9640 3460
rect 9864 3408 9916 3460
rect 10508 3476 10560 3528
rect 12532 3408 12584 3460
rect 6736 3340 6788 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 9772 3340 9824 3392
rect 11336 3340 11388 3392
rect 23664 3680 23716 3732
rect 24768 3680 24820 3732
rect 24860 3680 24912 3732
rect 13360 3612 13412 3664
rect 13636 3655 13688 3664
rect 13636 3621 13645 3655
rect 13645 3621 13679 3655
rect 13679 3621 13688 3655
rect 13636 3612 13688 3621
rect 14188 3612 14240 3664
rect 15660 3612 15712 3664
rect 15016 3544 15068 3596
rect 14556 3476 14608 3528
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 16764 3544 16816 3596
rect 19524 3544 19576 3596
rect 24860 3544 24912 3596
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 22284 3476 22336 3528
rect 23020 3476 23072 3528
rect 24676 3476 24728 3528
rect 24952 3476 25004 3528
rect 16120 3408 16172 3460
rect 17408 3408 17460 3460
rect 25964 3476 26016 3528
rect 12716 3383 12768 3392
rect 12716 3349 12725 3383
rect 12725 3349 12759 3383
rect 12759 3349 12768 3383
rect 12716 3340 12768 3349
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 13912 3340 13964 3392
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 21548 3340 21600 3392
rect 22836 3340 22888 3392
rect 25872 3408 25924 3460
rect 4703 3238 4755 3290
rect 4767 3238 4819 3290
rect 4831 3238 4883 3290
rect 4895 3238 4947 3290
rect 4959 3238 5011 3290
rect 10890 3238 10942 3290
rect 10954 3238 11006 3290
rect 11018 3238 11070 3290
rect 11082 3238 11134 3290
rect 11146 3238 11198 3290
rect 17077 3238 17129 3290
rect 17141 3238 17193 3290
rect 17205 3238 17257 3290
rect 17269 3238 17321 3290
rect 17333 3238 17385 3290
rect 23264 3238 23316 3290
rect 23328 3238 23380 3290
rect 23392 3238 23444 3290
rect 23456 3238 23508 3290
rect 23520 3238 23572 3290
rect 3056 3136 3108 3188
rect 4528 3136 4580 3188
rect 6000 3136 6052 3188
rect 6828 3136 6880 3188
rect 7104 3136 7156 3188
rect 7288 3136 7340 3188
rect 8300 3136 8352 3188
rect 8944 3136 8996 3188
rect 2596 3111 2648 3120
rect 2596 3077 2605 3111
rect 2605 3077 2639 3111
rect 2639 3077 2648 3111
rect 2596 3068 2648 3077
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2780 3000 2832 3052
rect 664 2932 716 2984
rect 5816 2932 5868 2984
rect 1952 2864 2004 2916
rect 20 2796 72 2848
rect 5448 2864 5500 2916
rect 6552 2864 6604 2916
rect 7748 3000 7800 3052
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 9772 3068 9824 3120
rect 10048 3136 10100 3188
rect 10784 3136 10836 3188
rect 12164 3136 12216 3188
rect 10508 3068 10560 3120
rect 11796 3111 11848 3120
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 9588 3000 9640 3052
rect 9312 2932 9364 2984
rect 9772 2932 9824 2984
rect 11244 3000 11296 3052
rect 11520 2864 11572 2916
rect 13268 3136 13320 3188
rect 14280 3136 14332 3188
rect 15568 3136 15620 3188
rect 17408 3136 17460 3188
rect 20904 3179 20956 3188
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 22008 3136 22060 3188
rect 14096 3068 14148 3120
rect 14924 3068 14976 3120
rect 17684 3068 17736 3120
rect 22100 3068 22152 3120
rect 22836 3068 22888 3120
rect 23112 3068 23164 3120
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 15476 2932 15528 2984
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 21732 3000 21784 3052
rect 20996 2932 21048 2984
rect 17040 2907 17092 2916
rect 17040 2873 17049 2907
rect 17049 2873 17083 2907
rect 17083 2873 17092 2907
rect 17040 2864 17092 2873
rect 17500 2864 17552 2916
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 24676 3000 24728 3052
rect 24676 2864 24728 2916
rect 9404 2796 9456 2848
rect 11336 2796 11388 2848
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 15384 2796 15436 2848
rect 16856 2796 16908 2848
rect 25136 2796 25188 2848
rect 4043 2694 4095 2746
rect 4107 2694 4159 2746
rect 4171 2694 4223 2746
rect 4235 2694 4287 2746
rect 4299 2694 4351 2746
rect 10230 2694 10282 2746
rect 10294 2694 10346 2746
rect 10358 2694 10410 2746
rect 10422 2694 10474 2746
rect 10486 2694 10538 2746
rect 16417 2694 16469 2746
rect 16481 2694 16533 2746
rect 16545 2694 16597 2746
rect 16609 2694 16661 2746
rect 16673 2694 16725 2746
rect 22604 2694 22656 2746
rect 22668 2694 22720 2746
rect 22732 2694 22784 2746
rect 22796 2694 22848 2746
rect 22860 2694 22912 2746
rect 1308 2592 1360 2644
rect 5172 2592 5224 2644
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 10784 2592 10836 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 12808 2592 12860 2644
rect 13820 2592 13872 2644
rect 15108 2592 15160 2644
rect 17040 2592 17092 2644
rect 21272 2592 21324 2644
rect 21916 2592 21968 2644
rect 1308 2320 1360 2372
rect 5448 2456 5500 2508
rect 12440 2456 12492 2508
rect 4068 2388 4120 2440
rect 6460 2388 6512 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 9036 2388 9088 2440
rect 10140 2388 10192 2440
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 12256 2431 12308 2440
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 13912 2524 13964 2576
rect 15936 2456 15988 2508
rect 17776 2524 17828 2576
rect 18972 2524 19024 2576
rect 20352 2524 20404 2576
rect 17684 2456 17736 2508
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 15384 2388 15436 2440
rect 15476 2388 15528 2440
rect 3884 2363 3936 2372
rect 3884 2329 3893 2363
rect 3893 2329 3927 2363
rect 3927 2329 3936 2363
rect 3884 2320 3936 2329
rect 5172 2320 5224 2372
rect 5356 2363 5408 2372
rect 5356 2329 5365 2363
rect 5365 2329 5399 2363
rect 5399 2329 5408 2363
rect 5356 2320 5408 2329
rect 3424 2252 3476 2304
rect 4620 2252 4672 2304
rect 5264 2252 5316 2304
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 9680 2252 9732 2304
rect 15660 2320 15712 2372
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 16856 2388 16908 2440
rect 19524 2388 19576 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 19340 2363 19392 2372
rect 19340 2329 19349 2363
rect 19349 2329 19383 2363
rect 19383 2329 19392 2363
rect 19340 2320 19392 2329
rect 20444 2388 20496 2440
rect 21732 2388 21784 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 22928 2431 22980 2440
rect 22928 2397 22937 2431
rect 22937 2397 22971 2431
rect 22971 2397 22980 2431
rect 22928 2388 22980 2397
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 24860 2388 24912 2440
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 12900 2252 12952 2304
rect 14924 2252 14976 2304
rect 15476 2252 15528 2304
rect 16488 2252 16540 2304
rect 18052 2252 18104 2304
rect 18788 2252 18840 2304
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 21732 2252 21784 2304
rect 24860 2295 24912 2304
rect 24860 2261 24869 2295
rect 24869 2261 24903 2295
rect 24903 2261 24912 2295
rect 24860 2252 24912 2261
rect 25228 2295 25280 2304
rect 25228 2261 25237 2295
rect 25237 2261 25271 2295
rect 25271 2261 25280 2295
rect 25228 2252 25280 2261
rect 4703 2150 4755 2202
rect 4767 2150 4819 2202
rect 4831 2150 4883 2202
rect 4895 2150 4947 2202
rect 4959 2150 5011 2202
rect 10890 2150 10942 2202
rect 10954 2150 11006 2202
rect 11018 2150 11070 2202
rect 11082 2150 11134 2202
rect 11146 2150 11198 2202
rect 17077 2150 17129 2202
rect 17141 2150 17193 2202
rect 17205 2150 17257 2202
rect 17269 2150 17321 2202
rect 17333 2150 17385 2202
rect 23264 2150 23316 2202
rect 23328 2150 23380 2202
rect 23392 2150 23444 2202
rect 23456 2150 23508 2202
rect 23520 2150 23572 2202
rect 5172 2048 5224 2100
rect 5356 1980 5408 2032
rect 5448 1980 5500 2032
rect 7380 2048 7432 2100
rect 12716 1980 12768 2032
rect 22928 2048 22980 2100
rect 8116 1912 8168 1964
rect 22376 1980 22428 2032
rect 19984 1912 20036 1964
rect 12624 1844 12676 1896
rect 12992 1844 13044 1896
rect 19340 1844 19392 1896
rect 13452 1776 13504 1828
rect 12440 1640 12492 1692
rect 22468 1640 22520 1692
rect 13268 1504 13320 1556
rect 24584 1504 24636 1556
rect 25780 1504 25832 1556
<< metal2 >>
rect 18 28381 74 29181
rect 662 28381 718 29181
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 32 25702 60 28381
rect 676 25974 704 28381
rect 1398 27024 1454 27033
rect 1398 26959 1454 26968
rect 1032 26036 1084 26042
rect 1032 25978 1084 25984
rect 664 25968 716 25974
rect 1044 25945 1072 25978
rect 664 25910 716 25916
rect 1030 25936 1086 25945
rect 1030 25871 1086 25880
rect 20 25696 72 25702
rect 20 25638 72 25644
rect 1412 25498 1440 26959
rect 1596 26586 1624 28591
rect 1950 28506 2006 29181
rect 2594 28506 2650 29181
rect 1950 28478 2268 28506
rect 1950 28381 2006 28478
rect 2240 26586 2268 28478
rect 2594 28478 2728 28506
rect 2594 28381 2650 28478
rect 1584 26580 1636 26586
rect 1584 26522 1636 26528
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2700 26450 2728 28478
rect 3238 28381 3294 29181
rect 3882 28381 3938 29181
rect 5170 28381 5226 29181
rect 5814 28381 5870 29181
rect 6458 28381 6514 29181
rect 7102 28506 7158 29181
rect 7102 28478 7420 28506
rect 7102 28381 7158 28478
rect 2870 26616 2926 26625
rect 2870 26551 2926 26560
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 1768 26308 1820 26314
rect 1768 26250 1820 26256
rect 1400 25492 1452 25498
rect 1400 25434 1452 25440
rect 1032 25288 1084 25294
rect 1030 25256 1032 25265
rect 1084 25256 1086 25265
rect 1030 25191 1086 25200
rect 940 24132 992 24138
rect 940 24074 992 24080
rect 952 23905 980 24074
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 938 23896 994 23905
rect 1596 23866 1624 24006
rect 938 23831 994 23840
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23497 1440 23666
rect 1582 23624 1638 23633
rect 1582 23559 1584 23568
rect 1636 23559 1638 23568
rect 1584 23530 1636 23536
rect 1398 23488 1454 23497
rect 1398 23423 1454 23432
rect 938 22536 994 22545
rect 938 22471 994 22480
rect 952 22438 980 22471
rect 940 22432 992 22438
rect 940 22374 992 22380
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 952 21185 980 21286
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20641 1440 20878
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 1596 19666 1624 20742
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1412 19638 1624 19666
rect 1412 18170 1440 19638
rect 1582 19544 1638 19553
rect 1582 19479 1584 19488
rect 1636 19479 1638 19488
rect 1584 19450 1636 19456
rect 1490 19408 1546 19417
rect 1490 19343 1492 19352
rect 1544 19343 1546 19352
rect 1492 19314 1544 19320
rect 1490 18320 1546 18329
rect 1490 18255 1492 18264
rect 1544 18255 1546 18264
rect 1492 18226 1544 18232
rect 1412 18142 1532 18170
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 940 17128 992 17134
rect 938 17096 940 17105
rect 992 17096 994 17105
rect 938 17031 994 17040
rect 1412 16561 1440 17138
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15745 980 15846
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 940 14408 992 14414
rect 938 14376 940 14385
rect 992 14376 994 14385
rect 938 14311 994 14320
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 952 13025 980 13126
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 1504 12434 1532 18142
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17921 1624 18022
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1688 17746 1716 19858
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1582 17096 1638 17105
rect 1582 17031 1584 17040
rect 1636 17031 1638 17040
rect 1584 17002 1636 17008
rect 1688 16794 1716 17682
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 15162 1716 16730
rect 1780 15473 1808 26250
rect 2884 25906 2912 26551
rect 3252 26382 3280 28381
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 1872 19242 1900 25842
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3332 25696 3384 25702
rect 3332 25638 3384 25644
rect 2044 25220 2096 25226
rect 2044 25162 2096 25168
rect 2056 19904 2084 25162
rect 2688 25152 2740 25158
rect 2688 25094 2740 25100
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22234 2268 22374
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2136 21956 2188 21962
rect 2136 21898 2188 21904
rect 2148 21690 2176 21898
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2424 21690 2452 21830
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2332 21146 2360 21490
rect 2410 21448 2466 21457
rect 2410 21383 2466 21392
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2056 19876 2268 19904
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 2056 19514 2084 19722
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1964 19281 1992 19314
rect 1950 19272 2006 19281
rect 1860 19236 1912 19242
rect 1950 19207 2006 19216
rect 1860 19178 1912 19184
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2056 17746 2084 18022
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 1872 16153 1900 16934
rect 1858 16144 1914 16153
rect 1858 16079 1914 16088
rect 2056 15502 2084 16934
rect 2044 15496 2096 15502
rect 1766 15464 1822 15473
rect 2044 15438 2096 15444
rect 1766 15399 1822 15408
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1872 14618 1900 14894
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1504 12406 1716 12434
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 1412 11626 1440 12174
rect 938 11591 994 11600
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10305 980 10406
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 1412 10130 1440 11562
rect 1584 11008 1636 11014
rect 1582 10976 1584 10985
rect 1636 10976 1638 10985
rect 1582 10911 1638 10920
rect 1490 10704 1546 10713
rect 1490 10639 1492 10648
rect 1544 10639 1546 10648
rect 1492 10610 1544 10616
rect 1688 10169 1716 12406
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1872 10606 1900 11630
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1674 10160 1730 10169
rect 1400 10124 1452 10130
rect 1674 10095 1730 10104
rect 1400 10066 1452 10072
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 952 9382 980 9551
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 8265 1716 8298
rect 1674 8256 1730 8265
rect 1674 8191 1730 8200
rect 938 7576 994 7585
rect 938 7511 940 7520
rect 992 7511 994 7520
rect 940 7482 992 7488
rect 1872 7324 1900 10542
rect 2056 8498 2084 15438
rect 2148 12714 2176 19110
rect 2240 18154 2268 19876
rect 2424 18986 2452 21383
rect 2516 19394 2544 22578
rect 2700 20505 2728 25094
rect 3068 22778 3096 25638
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3344 22094 3372 25638
rect 3160 22066 3372 22094
rect 2964 20868 3016 20874
rect 2964 20810 3016 20816
rect 2686 20496 2742 20505
rect 2686 20431 2742 20440
rect 2976 20398 3004 20810
rect 2964 20392 3016 20398
rect 2962 20360 2964 20369
rect 3016 20360 3018 20369
rect 2962 20295 3018 20304
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2608 19514 2636 19994
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2700 19514 2728 19858
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2516 19366 2728 19394
rect 2424 18958 2636 18986
rect 2228 18148 2280 18154
rect 2228 18090 2280 18096
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2240 17338 2268 17546
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 14618 2452 14758
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2516 14414 2544 15982
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2424 11898 2452 12786
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10033 2176 11018
rect 2332 10538 2360 11562
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2134 10024 2190 10033
rect 2134 9959 2190 9968
rect 2332 9602 2360 10474
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 9994 2452 10406
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2332 9574 2452 9602
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7818 1992 8230
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 2056 7478 2084 8434
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2044 7336 2096 7342
rect 1872 7296 2044 7324
rect 2044 7278 2096 7284
rect 2056 6730 2084 7278
rect 2424 7274 2452 9574
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2516 7546 2544 8434
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2424 6866 2452 7210
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4865 980 5170
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 1582 4584 1638 4593
rect 952 4185 980 4558
rect 1582 4519 1638 4528
rect 1596 4486 1624 4519
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1032 3528 1084 3534
rect 1030 3496 1032 3505
rect 1084 3496 1086 3505
rect 1030 3431 1086 3440
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 676 800 704 2926
rect 1308 2644 1360 2650
rect 1308 2586 1360 2592
rect 1320 2530 1348 2586
rect 1228 2502 1348 2530
rect 1228 1170 1256 2502
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 1465 1348 2314
rect 1596 2145 1624 3334
rect 2608 3126 2636 18958
rect 2700 6254 2728 19366
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17338 2912 17478
rect 3068 17338 3096 18226
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3160 17218 3188 22066
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 3344 21146 3372 21558
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3252 20534 3280 21082
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 3252 20330 3280 20470
rect 3436 20346 3464 26250
rect 3608 23248 3660 23254
rect 3608 23190 3660 23196
rect 3620 22574 3648 23190
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3620 22234 3648 22510
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 3344 20318 3464 20346
rect 3344 19802 3372 20318
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3344 19774 3464 19802
rect 2780 17196 2832 17202
rect 3160 17190 3280 17218
rect 2780 17138 2832 17144
rect 2792 16182 2820 17138
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2884 15978 2912 16730
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 15162 2820 15302
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2884 14550 2912 15914
rect 3068 15502 3096 15982
rect 3160 15978 3188 17070
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3160 15026 3188 15914
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 2976 14618 3004 14962
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3068 14074 3096 14418
rect 3252 14278 3280 17190
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3344 14890 3372 15438
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3252 14074 3280 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2884 12986 2912 13670
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12374 2820 12718
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2884 12434 2912 12582
rect 3068 12442 3096 13194
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3056 12436 3108 12442
rect 2884 12406 3004 12434
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2792 11694 2820 12310
rect 2976 12170 3004 12406
rect 3056 12378 3108 12384
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 3160 12050 3188 13126
rect 3240 12436 3292 12442
rect 3436 12434 3464 19774
rect 3528 19446 3556 20198
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3620 19310 3648 20198
rect 3712 19922 3740 22714
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3804 22234 3832 22646
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3792 20460 3844 20466
rect 3792 20402 3844 20408
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3804 18970 3832 20402
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3528 16794 3556 17002
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3620 16674 3648 18770
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3712 17338 3740 17682
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3528 16646 3648 16674
rect 3528 15570 3556 16646
rect 3712 16590 3740 17002
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3620 16250 3648 16526
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3804 15638 3832 16458
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 15094 3556 15302
rect 3896 15094 3924 28381
rect 4043 26684 4351 26693
rect 4043 26682 4049 26684
rect 4105 26682 4129 26684
rect 4185 26682 4209 26684
rect 4265 26682 4289 26684
rect 4345 26682 4351 26684
rect 4105 26630 4107 26682
rect 4287 26630 4289 26682
rect 4043 26628 4049 26630
rect 4105 26628 4129 26630
rect 4185 26628 4209 26630
rect 4265 26628 4289 26630
rect 4345 26628 4351 26630
rect 4043 26619 4351 26628
rect 5184 26382 5212 28381
rect 5828 26382 5856 28381
rect 5908 26512 5960 26518
rect 5908 26454 5960 26460
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 4703 26140 5011 26149
rect 4703 26138 4709 26140
rect 4765 26138 4789 26140
rect 4845 26138 4869 26140
rect 4925 26138 4949 26140
rect 5005 26138 5011 26140
rect 4765 26086 4767 26138
rect 4947 26086 4949 26138
rect 4703 26084 4709 26086
rect 4765 26084 4789 26086
rect 4845 26084 4869 26086
rect 4925 26084 4949 26086
rect 5005 26084 5011 26086
rect 4703 26075 5011 26084
rect 4043 25596 4351 25605
rect 4043 25594 4049 25596
rect 4105 25594 4129 25596
rect 4185 25594 4209 25596
rect 4265 25594 4289 25596
rect 4345 25594 4351 25596
rect 4105 25542 4107 25594
rect 4287 25542 4289 25594
rect 4043 25540 4049 25542
rect 4105 25540 4129 25542
rect 4185 25540 4209 25542
rect 4265 25540 4289 25542
rect 4345 25540 4351 25542
rect 4043 25531 4351 25540
rect 4703 25052 5011 25061
rect 4703 25050 4709 25052
rect 4765 25050 4789 25052
rect 4845 25050 4869 25052
rect 4925 25050 4949 25052
rect 5005 25050 5011 25052
rect 4765 24998 4767 25050
rect 4947 24998 4949 25050
rect 4703 24996 4709 24998
rect 4765 24996 4789 24998
rect 4845 24996 4869 24998
rect 4925 24996 4949 24998
rect 5005 24996 5011 24998
rect 4703 24987 5011 24996
rect 4043 24508 4351 24517
rect 4043 24506 4049 24508
rect 4105 24506 4129 24508
rect 4185 24506 4209 24508
rect 4265 24506 4289 24508
rect 4345 24506 4351 24508
rect 4105 24454 4107 24506
rect 4287 24454 4289 24506
rect 4043 24452 4049 24454
rect 4105 24452 4129 24454
rect 4185 24452 4209 24454
rect 4265 24452 4289 24454
rect 4345 24452 4351 24454
rect 4043 24443 4351 24452
rect 4703 23964 5011 23973
rect 4703 23962 4709 23964
rect 4765 23962 4789 23964
rect 4845 23962 4869 23964
rect 4925 23962 4949 23964
rect 5005 23962 5011 23964
rect 4765 23910 4767 23962
rect 4947 23910 4949 23962
rect 4703 23908 4709 23910
rect 4765 23908 4789 23910
rect 4845 23908 4869 23910
rect 4925 23908 4949 23910
rect 5005 23908 5011 23910
rect 4703 23899 5011 23908
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 4043 23420 4351 23429
rect 4043 23418 4049 23420
rect 4105 23418 4129 23420
rect 4185 23418 4209 23420
rect 4265 23418 4289 23420
rect 4345 23418 4351 23420
rect 4105 23366 4107 23418
rect 4287 23366 4289 23418
rect 4043 23364 4049 23366
rect 4105 23364 4129 23366
rect 4185 23364 4209 23366
rect 4265 23364 4289 23366
rect 4345 23364 4351 23366
rect 4043 23355 4351 23364
rect 5276 22982 5304 23666
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4043 22332 4351 22341
rect 4043 22330 4049 22332
rect 4105 22330 4129 22332
rect 4185 22330 4209 22332
rect 4265 22330 4289 22332
rect 4345 22330 4351 22332
rect 4105 22278 4107 22330
rect 4287 22278 4289 22330
rect 4043 22276 4049 22278
rect 4105 22276 4129 22278
rect 4185 22276 4209 22278
rect 4265 22276 4289 22278
rect 4345 22276 4351 22278
rect 4043 22267 4351 22276
rect 4448 22234 4476 22442
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4043 21244 4351 21253
rect 4043 21242 4049 21244
rect 4105 21242 4129 21244
rect 4185 21242 4209 21244
rect 4265 21242 4289 21244
rect 4345 21242 4351 21244
rect 4105 21190 4107 21242
rect 4287 21190 4289 21242
rect 4043 21188 4049 21190
rect 4105 21188 4129 21190
rect 4185 21188 4209 21190
rect 4265 21188 4289 21190
rect 4345 21188 4351 21190
rect 4043 21179 4351 21188
rect 4448 21010 4476 21898
rect 4540 21622 4568 22374
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 4632 21554 4660 22918
rect 4703 22876 5011 22885
rect 4703 22874 4709 22876
rect 4765 22874 4789 22876
rect 4845 22874 4869 22876
rect 4925 22874 4949 22876
rect 5005 22874 5011 22876
rect 4765 22822 4767 22874
rect 4947 22822 4949 22874
rect 4703 22820 4709 22822
rect 4765 22820 4789 22822
rect 4845 22820 4869 22822
rect 4925 22820 4949 22822
rect 5005 22820 5011 22822
rect 4703 22811 5011 22820
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 4703 21788 5011 21797
rect 4703 21786 4709 21788
rect 4765 21786 4789 21788
rect 4845 21786 4869 21788
rect 4925 21786 4949 21788
rect 5005 21786 5011 21788
rect 4765 21734 4767 21786
rect 4947 21734 4949 21786
rect 4703 21732 4709 21734
rect 4765 21732 4789 21734
rect 4845 21732 4869 21734
rect 4925 21732 4949 21734
rect 5005 21732 5011 21734
rect 4703 21723 5011 21732
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4043 20156 4351 20165
rect 4043 20154 4049 20156
rect 4105 20154 4129 20156
rect 4185 20154 4209 20156
rect 4265 20154 4289 20156
rect 4345 20154 4351 20156
rect 4105 20102 4107 20154
rect 4287 20102 4289 20154
rect 4043 20100 4049 20102
rect 4105 20100 4129 20102
rect 4185 20100 4209 20102
rect 4265 20100 4289 20102
rect 4345 20100 4351 20102
rect 4043 20091 4351 20100
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4080 19922 4108 19994
rect 4250 19952 4306 19961
rect 4068 19916 4120 19922
rect 4250 19887 4252 19896
rect 4068 19858 4120 19864
rect 4304 19887 4306 19896
rect 4252 19858 4304 19864
rect 4448 19854 4476 20946
rect 5000 20874 5028 21286
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4703 20700 5011 20709
rect 4703 20698 4709 20700
rect 4765 20698 4789 20700
rect 4845 20698 4869 20700
rect 4925 20698 4949 20700
rect 5005 20698 5011 20700
rect 4765 20646 4767 20698
rect 4947 20646 4949 20698
rect 4703 20644 4709 20646
rect 4765 20644 4789 20646
rect 4845 20644 4869 20646
rect 4925 20644 4949 20646
rect 5005 20644 5011 20646
rect 4703 20635 5011 20644
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4528 19848 4580 19854
rect 4724 19802 4752 19994
rect 4816 19922 4844 20538
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 5092 19854 5120 22578
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 5184 21486 5212 21898
rect 5276 21554 5304 22918
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5184 20942 5212 21422
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 4528 19790 4580 19796
rect 4344 19780 4396 19786
rect 4344 19722 4396 19728
rect 4356 19514 4384 19722
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4540 19446 4568 19790
rect 4632 19774 4752 19802
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 4436 19440 4488 19446
rect 4436 19382 4488 19388
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4043 19068 4351 19077
rect 4043 19066 4049 19068
rect 4105 19066 4129 19068
rect 4185 19066 4209 19068
rect 4265 19066 4289 19068
rect 4345 19066 4351 19068
rect 4105 19014 4107 19066
rect 4287 19014 4289 19066
rect 4043 19012 4049 19014
rect 4105 19012 4129 19014
rect 4185 19012 4209 19014
rect 4265 19012 4289 19014
rect 4345 19012 4351 19014
rect 4043 19003 4351 19012
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4252 18896 4304 18902
rect 4158 18864 4214 18873
rect 4252 18838 4304 18844
rect 4158 18799 4214 18808
rect 4172 18698 4200 18799
rect 4264 18737 4292 18838
rect 4356 18834 4384 18906
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4250 18728 4306 18737
rect 4160 18692 4212 18698
rect 4250 18663 4306 18672
rect 4160 18634 4212 18640
rect 4344 18216 4396 18222
rect 4448 18204 4476 19382
rect 4528 19304 4580 19310
rect 4526 19272 4528 19281
rect 4580 19272 4582 19281
rect 4632 19242 4660 19774
rect 5276 19666 5304 20878
rect 5092 19638 5304 19666
rect 4703 19612 5011 19621
rect 4703 19610 4709 19612
rect 4765 19610 4789 19612
rect 4845 19610 4869 19612
rect 4925 19610 4949 19612
rect 5005 19610 5011 19612
rect 4765 19558 4767 19610
rect 4947 19558 4949 19610
rect 4703 19556 4709 19558
rect 4765 19556 4789 19558
rect 4845 19556 4869 19558
rect 4925 19556 4949 19558
rect 5005 19556 5011 19558
rect 4703 19547 5011 19556
rect 5092 19496 5120 19638
rect 5368 19496 5396 22102
rect 5460 19802 5488 26182
rect 5920 26042 5948 26454
rect 6472 26382 6500 28381
rect 7392 26586 7420 28478
rect 8390 28381 8446 29181
rect 9034 28506 9090 29181
rect 9034 28478 9352 28506
rect 9034 28381 9090 28478
rect 8404 26586 8432 28381
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 9324 26382 9352 28478
rect 9678 28381 9734 29181
rect 10966 28381 11022 29181
rect 11610 28381 11666 29181
rect 12254 28381 12310 29181
rect 12898 28381 12954 29181
rect 14186 28506 14242 29181
rect 14186 28478 14504 28506
rect 14186 28381 14242 28478
rect 9692 26382 9720 28381
rect 10980 27418 11008 28381
rect 10980 27390 11100 27418
rect 10230 26684 10538 26693
rect 10230 26682 10236 26684
rect 10292 26682 10316 26684
rect 10372 26682 10396 26684
rect 10452 26682 10476 26684
rect 10532 26682 10538 26684
rect 10292 26630 10294 26682
rect 10474 26630 10476 26682
rect 10230 26628 10236 26630
rect 10292 26628 10316 26630
rect 10372 26628 10396 26630
rect 10452 26628 10476 26630
rect 10532 26628 10538 26630
rect 10230 26619 10538 26628
rect 11072 26586 11100 27390
rect 11624 26586 11652 28381
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 10692 26512 10744 26518
rect 10692 26454 10744 26460
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 8208 26308 8260 26314
rect 8208 26250 8260 26256
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 6092 26240 6144 26246
rect 6736 26240 6788 26246
rect 6144 26200 6316 26228
rect 6092 26182 6144 26188
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23118 5580 23462
rect 5736 23118 5764 23598
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 5920 23118 5948 23530
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5552 22574 5580 23054
rect 5736 22778 5764 23054
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5736 21894 5764 22510
rect 5828 22234 5856 23054
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5644 21622 5672 21830
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5644 21468 5672 21558
rect 5724 21480 5776 21486
rect 5644 21440 5724 21468
rect 5724 21422 5776 21428
rect 5828 21418 5856 21966
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5552 21146 5580 21354
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5552 20942 5580 21082
rect 5920 21078 5948 21830
rect 6012 21622 6040 23598
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6000 21616 6052 21622
rect 6000 21558 6052 21564
rect 6104 21554 6132 23054
rect 6196 23050 6224 23666
rect 6184 23044 6236 23050
rect 6184 22986 6236 22992
rect 6196 22574 6224 22986
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5460 19774 5580 19802
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5000 19468 5120 19496
rect 5184 19468 5396 19496
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4526 19207 4582 19216
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18426 4568 19110
rect 4632 18766 4660 19178
rect 4816 19009 4844 19314
rect 4802 19000 4858 19009
rect 4802 18935 4858 18944
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4802 18864 4858 18873
rect 4724 18822 4802 18850
rect 4724 18766 4752 18822
rect 4802 18799 4858 18808
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4908 18630 4936 18906
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4896 18624 4948 18630
rect 5000 18612 5028 19468
rect 5184 19394 5212 19468
rect 5092 19366 5212 19394
rect 5264 19372 5316 19378
rect 5092 18970 5120 19366
rect 5264 19314 5316 19320
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5000 18584 5120 18612
rect 4896 18566 4948 18572
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4396 18176 4476 18204
rect 4344 18158 4396 18164
rect 4043 17980 4351 17989
rect 4043 17978 4049 17980
rect 4105 17978 4129 17980
rect 4185 17978 4209 17980
rect 4265 17978 4289 17980
rect 4345 17978 4351 17980
rect 4105 17926 4107 17978
rect 4287 17926 4289 17978
rect 4043 17924 4049 17926
rect 4105 17924 4129 17926
rect 4185 17924 4209 17926
rect 4265 17924 4289 17926
rect 4345 17924 4351 17926
rect 4043 17915 4351 17924
rect 4448 17882 4476 18176
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3988 16998 4016 17478
rect 4080 17202 4108 17614
rect 4448 17338 4476 17818
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4632 17270 4660 18566
rect 4703 18524 5011 18533
rect 4703 18522 4709 18524
rect 4765 18522 4789 18524
rect 4845 18522 4869 18524
rect 4925 18522 4949 18524
rect 5005 18522 5011 18524
rect 4765 18470 4767 18522
rect 4947 18470 4949 18522
rect 4703 18468 4709 18470
rect 4765 18468 4789 18470
rect 4845 18468 4869 18470
rect 4925 18468 4949 18470
rect 5005 18468 5011 18470
rect 4703 18459 5011 18468
rect 4703 17436 5011 17445
rect 4703 17434 4709 17436
rect 4765 17434 4789 17436
rect 4845 17434 4869 17436
rect 4925 17434 4949 17436
rect 5005 17434 5011 17436
rect 4765 17382 4767 17434
rect 4947 17382 4949 17434
rect 4703 17380 4709 17382
rect 4765 17380 4789 17382
rect 4845 17380 4869 17382
rect 4925 17380 4949 17382
rect 5005 17380 5011 17382
rect 4703 17371 5011 17380
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 4043 16892 4351 16901
rect 4043 16890 4049 16892
rect 4105 16890 4129 16892
rect 4185 16890 4209 16892
rect 4265 16890 4289 16892
rect 4345 16890 4351 16892
rect 4105 16838 4107 16890
rect 4287 16838 4289 16890
rect 4043 16836 4049 16838
rect 4105 16836 4129 16838
rect 4185 16836 4209 16838
rect 4265 16836 4289 16838
rect 4345 16836 4351 16838
rect 4043 16827 4351 16836
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16182 4108 16390
rect 4264 16250 4292 16662
rect 4540 16250 4568 16662
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4632 16182 4660 16458
rect 4703 16348 5011 16357
rect 4703 16346 4709 16348
rect 4765 16346 4789 16348
rect 4845 16346 4869 16348
rect 4925 16346 4949 16348
rect 5005 16346 5011 16348
rect 4765 16294 4767 16346
rect 4947 16294 4949 16346
rect 4703 16292 4709 16294
rect 4765 16292 4789 16294
rect 4845 16292 4869 16294
rect 4925 16292 4949 16294
rect 5005 16292 5011 16294
rect 4703 16283 5011 16292
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4043 15804 4351 15813
rect 4043 15802 4049 15804
rect 4105 15802 4129 15804
rect 4185 15802 4209 15804
rect 4265 15802 4289 15804
rect 4345 15802 4351 15804
rect 4105 15750 4107 15802
rect 4287 15750 4289 15802
rect 4043 15748 4049 15750
rect 4105 15748 4129 15750
rect 4185 15748 4209 15750
rect 4265 15748 4289 15750
rect 4345 15748 4351 15750
rect 4043 15739 4351 15748
rect 4703 15260 5011 15269
rect 4703 15258 4709 15260
rect 4765 15258 4789 15260
rect 4845 15258 4869 15260
rect 4925 15258 4949 15260
rect 5005 15258 5011 15260
rect 4765 15206 4767 15258
rect 4947 15206 4949 15258
rect 4703 15204 4709 15206
rect 4765 15204 4789 15206
rect 4845 15204 4869 15206
rect 4925 15204 4949 15206
rect 5005 15204 5011 15206
rect 4703 15195 5011 15204
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 3884 15088 3936 15094
rect 3884 15030 3936 15036
rect 5092 14822 5120 18584
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4043 14716 4351 14725
rect 4043 14714 4049 14716
rect 4105 14714 4129 14716
rect 4185 14714 4209 14716
rect 4265 14714 4289 14716
rect 4345 14714 4351 14716
rect 4105 14662 4107 14714
rect 4287 14662 4289 14714
rect 4043 14660 4049 14662
rect 4105 14660 4129 14662
rect 4185 14660 4209 14662
rect 4265 14660 4289 14662
rect 4345 14660 4351 14662
rect 4043 14651 4351 14660
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13394 3832 13806
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3436 12406 3648 12434
rect 3240 12378 3292 12384
rect 3068 12022 3188 12050
rect 3068 11830 3096 12022
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 3252 11218 3280 12378
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10266 3556 10406
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9518 3188 9862
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3344 9178 3372 9454
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8430 3464 8910
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 7886 2820 8298
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7954 3556 8230
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3620 7750 3648 12406
rect 3896 12306 3924 14350
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4043 13628 4351 13637
rect 4043 13626 4049 13628
rect 4105 13626 4129 13628
rect 4185 13626 4209 13628
rect 4265 13626 4289 13628
rect 4345 13626 4351 13628
rect 4105 13574 4107 13626
rect 4287 13574 4289 13626
rect 4043 13572 4049 13574
rect 4105 13572 4129 13574
rect 4185 13572 4209 13574
rect 4265 13572 4289 13574
rect 4345 13572 4351 13574
rect 4043 13563 4351 13572
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4356 13297 4384 13330
rect 4342 13288 4398 13297
rect 4342 13223 4398 13232
rect 4448 12986 4476 13874
rect 4540 13326 4568 14282
rect 4632 14074 4660 14758
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4703 14172 5011 14181
rect 4703 14170 4709 14172
rect 4765 14170 4789 14172
rect 4845 14170 4869 14172
rect 4925 14170 4949 14172
rect 5005 14170 5011 14172
rect 4765 14118 4767 14170
rect 4947 14118 4949 14170
rect 4703 14116 4709 14118
rect 4765 14116 4789 14118
rect 4845 14116 4869 14118
rect 4925 14116 4949 14118
rect 5005 14116 5011 14118
rect 4703 14107 5011 14116
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 5092 13870 5120 14282
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13394 5120 13806
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 5184 13190 5212 19110
rect 5276 18902 5304 19314
rect 5368 18970 5396 19314
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5264 18896 5316 18902
rect 5262 18864 5264 18873
rect 5316 18864 5318 18873
rect 5262 18799 5318 18808
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5262 17912 5318 17921
rect 5262 17847 5318 17856
rect 5276 17678 5304 17847
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5368 17490 5396 18634
rect 5460 17785 5488 19654
rect 5446 17776 5502 17785
rect 5446 17711 5502 17720
rect 5552 17649 5580 19774
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 18902 5856 19110
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5538 17640 5594 17649
rect 5538 17575 5594 17584
rect 5276 17462 5396 17490
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4043 12540 4351 12549
rect 4043 12538 4049 12540
rect 4105 12538 4129 12540
rect 4185 12538 4209 12540
rect 4265 12538 4289 12540
rect 4345 12538 4351 12540
rect 4105 12486 4107 12538
rect 4287 12486 4289 12538
rect 4043 12484 4049 12486
rect 4105 12484 4129 12486
rect 4185 12484 4209 12486
rect 4265 12484 4289 12486
rect 4345 12484 4351 12486
rect 4043 12475 4351 12484
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 4540 11898 4568 13126
rect 4632 12918 4660 13126
rect 4703 13084 5011 13093
rect 4703 13082 4709 13084
rect 4765 13082 4789 13084
rect 4845 13082 4869 13084
rect 4925 13082 4949 13084
rect 5005 13082 5011 13084
rect 4765 13030 4767 13082
rect 4947 13030 4949 13082
rect 4703 13028 4709 13030
rect 4765 13028 4789 13030
rect 4845 13028 4869 13030
rect 4925 13028 4949 13030
rect 5005 13028 5011 13030
rect 4703 13019 5011 13028
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4724 12730 4752 12922
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4632 12702 4752 12730
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4043 11452 4351 11461
rect 4043 11450 4049 11452
rect 4105 11450 4129 11452
rect 4185 11450 4209 11452
rect 4265 11450 4289 11452
rect 4345 11450 4351 11452
rect 4105 11398 4107 11450
rect 4287 11398 4289 11450
rect 4043 11396 4049 11398
rect 4105 11396 4129 11398
rect 4185 11396 4209 11398
rect 4265 11396 4289 11398
rect 4345 11396 4351 11398
rect 4043 11387 4351 11396
rect 4540 11354 4568 11834
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4540 11150 4568 11290
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10674 4200 11018
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4043 10364 4351 10373
rect 4043 10362 4049 10364
rect 4105 10362 4129 10364
rect 4185 10362 4209 10364
rect 4265 10362 4289 10364
rect 4345 10362 4351 10364
rect 4105 10310 4107 10362
rect 4287 10310 4289 10362
rect 4043 10308 4049 10310
rect 4105 10308 4129 10310
rect 4185 10308 4209 10310
rect 4265 10308 4289 10310
rect 4345 10308 4351 10310
rect 4043 10299 4351 10308
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9586 3924 9862
rect 4632 9674 4660 12702
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12306 4752 12582
rect 4908 12442 4936 12786
rect 5092 12782 5120 13126
rect 5276 13002 5304 17462
rect 5736 17066 5764 18702
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 16561 5488 16594
rect 5446 16552 5502 16561
rect 5446 16487 5448 16496
rect 5500 16487 5502 16496
rect 5448 16458 5500 16464
rect 5460 15026 5488 16458
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5552 14890 5580 16662
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5644 15570 5672 15846
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5736 15434 5764 15846
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5368 13870 5396 14486
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14006 5580 14350
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5368 13326 5396 13670
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5184 12974 5304 13002
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4703 11996 5011 12005
rect 4703 11994 4709 11996
rect 4765 11994 4789 11996
rect 4845 11994 4869 11996
rect 4925 11994 4949 11996
rect 5005 11994 5011 11996
rect 4765 11942 4767 11994
rect 4947 11942 4949 11994
rect 4703 11940 4709 11942
rect 4765 11940 4789 11942
rect 4845 11940 4869 11942
rect 4925 11940 4949 11942
rect 5005 11940 5011 11942
rect 4703 11931 5011 11940
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5092 11626 5120 11834
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4703 10908 5011 10917
rect 4703 10906 4709 10908
rect 4765 10906 4789 10908
rect 4845 10906 4869 10908
rect 4925 10906 4949 10908
rect 5005 10906 5011 10908
rect 4765 10854 4767 10906
rect 4947 10854 4949 10906
rect 4703 10852 4709 10854
rect 4765 10852 4789 10854
rect 4845 10852 4869 10854
rect 4925 10852 4949 10854
rect 5005 10852 5011 10854
rect 4703 10843 5011 10852
rect 5092 10674 5120 10950
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 9926 4844 10542
rect 4908 10266 4936 10610
rect 5078 10568 5134 10577
rect 5078 10503 5134 10512
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4703 9820 5011 9829
rect 4703 9818 4709 9820
rect 4765 9818 4789 9820
rect 4845 9818 4869 9820
rect 4925 9818 4949 9820
rect 5005 9818 5011 9820
rect 4765 9766 4767 9818
rect 4947 9766 4949 9818
rect 4703 9764 4709 9766
rect 4765 9764 4789 9766
rect 4845 9764 4869 9766
rect 4925 9764 4949 9766
rect 5005 9764 5011 9766
rect 4703 9755 5011 9764
rect 4632 9654 4752 9674
rect 4632 9648 4764 9654
rect 4632 9646 4712 9648
rect 4250 9616 4306 9625
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 4160 9580 4212 9586
rect 4712 9590 4764 9596
rect 4250 9551 4252 9560
rect 4160 9522 4212 9528
rect 4304 9551 4306 9560
rect 4252 9522 4304 9528
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 8498 3740 9318
rect 3896 8974 3924 9522
rect 4172 9466 4200 9522
rect 4172 9438 4568 9466
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4043 9276 4351 9285
rect 4043 9274 4049 9276
rect 4105 9274 4129 9276
rect 4185 9274 4209 9276
rect 4265 9274 4289 9276
rect 4345 9274 4351 9276
rect 4105 9222 4107 9274
rect 4287 9222 4289 9274
rect 4043 9220 4049 9222
rect 4105 9220 4129 9222
rect 4185 9220 4209 9222
rect 4265 9220 4289 9222
rect 4345 9220 4351 9222
rect 4043 9211 4351 9220
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8634 3832 8774
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3896 8498 3924 8910
rect 4172 8498 4200 9046
rect 4448 9042 4476 9318
rect 4540 9042 4568 9438
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4356 8362 4384 8978
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8498 4476 8774
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4540 8242 4568 8978
rect 4632 8498 4660 9318
rect 4724 9110 4752 9590
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4703 8732 5011 8741
rect 4703 8730 4709 8732
rect 4765 8730 4789 8732
rect 4845 8730 4869 8732
rect 4925 8730 4949 8732
rect 5005 8730 5011 8732
rect 4765 8678 4767 8730
rect 4947 8678 4949 8730
rect 4703 8676 4709 8678
rect 4765 8676 4789 8678
rect 4845 8676 4869 8678
rect 4925 8676 4949 8678
rect 5005 8676 5011 8678
rect 4703 8667 5011 8676
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4540 8214 4660 8242
rect 4043 8188 4351 8197
rect 4043 8186 4049 8188
rect 4105 8186 4129 8188
rect 4185 8186 4209 8188
rect 4265 8186 4289 8188
rect 4345 8186 4351 8188
rect 4105 8134 4107 8186
rect 4287 8134 4289 8186
rect 4043 8132 4049 8134
rect 4105 8132 4129 8134
rect 4185 8132 4209 8134
rect 4265 8132 4289 8134
rect 4345 8132 4351 8134
rect 4043 8123 4351 8132
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 6905 2820 7346
rect 3068 7342 3096 7686
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 3068 3194 3096 7278
rect 3804 6798 3832 8026
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4043 7100 4351 7109
rect 4043 7098 4049 7100
rect 4105 7098 4129 7100
rect 4185 7098 4209 7100
rect 4265 7098 4289 7100
rect 4345 7098 4351 7100
rect 4105 7046 4107 7098
rect 4287 7046 4289 7098
rect 4043 7044 4049 7046
rect 4105 7044 4129 7046
rect 4185 7044 4209 7046
rect 4265 7044 4289 7046
rect 4345 7044 4351 7046
rect 4043 7035 4351 7044
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 4043 6012 4351 6021
rect 4043 6010 4049 6012
rect 4105 6010 4129 6012
rect 4185 6010 4209 6012
rect 4265 6010 4289 6012
rect 4345 6010 4351 6012
rect 4105 5958 4107 6010
rect 4287 5958 4289 6010
rect 4043 5956 4049 5958
rect 4105 5956 4129 5958
rect 4185 5956 4209 5958
rect 4265 5956 4289 5958
rect 4345 5956 4351 5958
rect 4043 5947 4351 5956
rect 4448 5710 4476 7958
rect 4632 7886 4660 8214
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4724 7818 4752 8366
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 7954 4844 8230
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4703 7644 5011 7653
rect 4703 7642 4709 7644
rect 4765 7642 4789 7644
rect 4845 7642 4869 7644
rect 4925 7642 4949 7644
rect 5005 7642 5011 7644
rect 4765 7590 4767 7642
rect 4947 7590 4949 7642
rect 4703 7588 4709 7590
rect 4765 7588 4789 7590
rect 4845 7588 4869 7590
rect 4925 7588 4949 7590
rect 5005 7588 5011 7590
rect 4703 7579 5011 7588
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 6746 4660 7142
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4540 6718 4660 6746
rect 4540 6322 4568 6718
rect 4724 6644 4752 6870
rect 4632 6616 4752 6644
rect 4528 6316 4580 6322
rect 4632 6304 4660 6616
rect 4703 6556 5011 6565
rect 4703 6554 4709 6556
rect 4765 6554 4789 6556
rect 4845 6554 4869 6556
rect 4925 6554 4949 6556
rect 5005 6554 5011 6556
rect 4765 6502 4767 6554
rect 4947 6502 4949 6554
rect 4703 6500 4709 6502
rect 4765 6500 4789 6502
rect 4845 6500 4869 6502
rect 4925 6500 4949 6502
rect 5005 6500 5011 6502
rect 4703 6491 5011 6500
rect 4712 6316 4764 6322
rect 4632 6276 4712 6304
rect 4528 6258 4580 6264
rect 4712 6258 4764 6264
rect 5092 6202 5120 10503
rect 4540 6174 5120 6202
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5370 4476 5646
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4043 4924 4351 4933
rect 4043 4922 4049 4924
rect 4105 4922 4129 4924
rect 4185 4922 4209 4924
rect 4265 4922 4289 4924
rect 4345 4922 4351 4924
rect 4105 4870 4107 4922
rect 4287 4870 4289 4922
rect 4043 4868 4049 4870
rect 4105 4868 4129 4870
rect 4185 4868 4209 4870
rect 4265 4868 4289 4870
rect 4345 4868 4351 4870
rect 4043 4859 4351 4868
rect 4043 3836 4351 3845
rect 4043 3834 4049 3836
rect 4105 3834 4129 3836
rect 4185 3834 4209 3836
rect 4265 3834 4289 3836
rect 4345 3834 4351 3836
rect 4105 3782 4107 3834
rect 4287 3782 4289 3834
rect 4043 3780 4049 3782
rect 4105 3780 4129 3782
rect 4185 3780 4209 3782
rect 4265 3780 4289 3782
rect 4345 3780 4351 3782
rect 4043 3771 4351 3780
rect 4448 3466 4476 5306
rect 4540 3618 4568 6174
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4632 5166 4660 6054
rect 4703 5468 5011 5477
rect 4703 5466 4709 5468
rect 4765 5466 4789 5468
rect 4845 5466 4869 5468
rect 4925 5466 4949 5468
rect 5005 5466 5011 5468
rect 4765 5414 4767 5466
rect 4947 5414 4949 5466
rect 4703 5412 4709 5414
rect 4765 5412 4789 5414
rect 4845 5412 4869 5414
rect 4925 5412 4949 5414
rect 5005 5412 5011 5414
rect 4703 5403 5011 5412
rect 5092 5370 5120 6054
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4703 4380 5011 4389
rect 4703 4378 4709 4380
rect 4765 4378 4789 4380
rect 4845 4378 4869 4380
rect 4925 4378 4949 4380
rect 5005 4378 5011 4380
rect 4765 4326 4767 4378
rect 4947 4326 4949 4378
rect 4703 4324 4709 4326
rect 4765 4324 4789 4326
rect 4845 4324 4869 4326
rect 4925 4324 4949 4326
rect 5005 4324 5011 4326
rect 4703 4315 5011 4324
rect 4540 3590 4660 3618
rect 4632 3466 4660 3590
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4540 3194 4568 3402
rect 4703 3292 5011 3301
rect 4703 3290 4709 3292
rect 4765 3290 4789 3292
rect 4845 3290 4869 3292
rect 4925 3290 4949 3292
rect 5005 3290 5011 3292
rect 4765 3238 4767 3290
rect 4947 3238 4949 3290
rect 4703 3236 4709 3238
rect 4765 3236 4789 3238
rect 4845 3236 4869 3238
rect 4925 3236 4949 3238
rect 5005 3236 5011 3238
rect 4703 3227 5011 3236
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 2596 3120 2648 3126
rect 2042 3088 2098 3097
rect 2596 3062 2648 3068
rect 2042 3023 2044 3032
rect 2096 3023 2098 3032
rect 2780 3052 2832 3058
rect 2044 2994 2096 3000
rect 2780 2994 2832 3000
rect 1952 2916 2004 2922
rect 1952 2858 2004 2864
rect 1582 2136 1638 2145
rect 1582 2071 1638 2080
rect 1306 1456 1362 1465
rect 1306 1391 1362 1400
rect 1228 1142 1348 1170
rect 1320 800 1348 1142
rect 1964 800 1992 2858
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2792 785 2820 2994
rect 4043 2748 4351 2757
rect 4043 2746 4049 2748
rect 4105 2746 4129 2748
rect 4185 2746 4209 2748
rect 4265 2746 4289 2748
rect 4345 2746 4351 2748
rect 4105 2694 4107 2746
rect 4287 2694 4289 2746
rect 4043 2692 4049 2694
rect 4105 2692 4129 2694
rect 4185 2692 4209 2694
rect 4265 2692 4289 2694
rect 4345 2692 4351 2694
rect 4043 2683 4351 2692
rect 5184 2650 5212 12974
rect 5368 12628 5396 13126
rect 5460 12696 5488 13670
rect 5460 12668 5580 12696
rect 5276 12600 5396 12628
rect 5276 6202 5304 12600
rect 5552 12238 5580 12668
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10674 5396 10950
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 10062 5396 10610
rect 5460 10266 5488 11086
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10742 5580 10950
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5538 10568 5594 10577
rect 5644 10554 5672 14758
rect 5828 12434 5856 18838
rect 5920 17338 5948 19382
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18086 6132 18702
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6012 16794 6040 17206
rect 6104 16998 6132 18022
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5920 15162 5948 16050
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 13938 6040 14214
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6196 13462 6224 13738
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6288 13410 6316 26200
rect 6564 26200 6736 26228
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6380 24954 6408 25230
rect 6368 24948 6420 24954
rect 6368 24890 6420 24896
rect 6368 23180 6420 23186
rect 6368 23122 6420 23128
rect 6380 21622 6408 23122
rect 6564 21978 6592 26200
rect 6736 26182 6788 26188
rect 6736 24880 6788 24886
rect 6840 24857 6868 26250
rect 6736 24822 6788 24828
rect 6826 24848 6882 24857
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6656 22778 6684 23122
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6472 21950 6592 21978
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6472 19802 6500 21950
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21554 6592 21830
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6564 21146 6592 21490
rect 6656 21486 6684 21966
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6656 20806 6684 21422
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6472 19774 6592 19802
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19514 6500 19654
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6380 16794 6408 18294
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14482 6408 14758
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 14074 6408 14282
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6564 13802 6592 19774
rect 6656 19378 6684 19994
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6656 17134 6684 18906
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6458 13424 6514 13433
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5736 12406 5856 12434
rect 5736 11218 5764 12406
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5594 10526 5672 10554
rect 5538 10503 5594 10512
rect 5632 10464 5684 10470
rect 5552 10424 5632 10452
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8634 5396 8978
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5356 6792 5408 6798
rect 5354 6760 5356 6769
rect 5408 6760 5410 6769
rect 5460 6746 5488 9658
rect 5552 9586 5580 10424
rect 5632 10406 5684 10412
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9586 5672 9930
rect 5736 9586 5764 10610
rect 5828 9625 5856 12038
rect 5920 11762 5948 13330
rect 6092 12232 6144 12238
rect 6090 12200 6092 12209
rect 6144 12200 6146 12209
rect 6090 12135 6146 12144
rect 6196 11898 6224 13398
rect 6288 13382 6458 13410
rect 6458 13359 6514 13368
rect 6748 12434 6776 24822
rect 6826 24783 6828 24792
rect 6880 24783 6882 24792
rect 6828 24754 6880 24760
rect 7300 24698 7328 26250
rect 8116 25832 8168 25838
rect 8116 25774 8168 25780
rect 8128 25430 8156 25774
rect 8220 25498 8248 26250
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 9036 25968 9088 25974
rect 9036 25910 9088 25916
rect 8300 25832 8352 25838
rect 8588 25809 8616 25910
rect 8668 25832 8720 25838
rect 8300 25774 8352 25780
rect 8574 25800 8630 25809
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 8116 25424 8168 25430
rect 8116 25366 8168 25372
rect 7656 24880 7708 24886
rect 7656 24822 7708 24828
rect 7300 24670 7512 24698
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 24410 7328 24550
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 23322 6868 23462
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 6840 22030 6868 22918
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6932 22234 6960 22510
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6826 20224 6882 20233
rect 6826 20159 6882 20168
rect 6840 19990 6868 20159
rect 6828 19984 6880 19990
rect 6828 19926 6880 19932
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 19378 6868 19722
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6920 19372 6972 19378
rect 7024 19360 7052 22646
rect 7116 21622 7144 22918
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7208 21622 7236 22578
rect 7300 22234 7328 22918
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7196 21616 7248 21622
rect 7196 21558 7248 21564
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7116 21078 7144 21422
rect 7300 21146 7328 21966
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7104 21072 7156 21078
rect 7104 21014 7156 21020
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19990 7144 20334
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19378 7144 19790
rect 7208 19446 7236 20198
rect 7300 20058 7328 21082
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 7286 19952 7342 19961
rect 7286 19887 7342 19896
rect 7300 19718 7328 19887
rect 7392 19854 7420 20742
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 6972 19332 7052 19360
rect 7104 19372 7156 19378
rect 6920 19314 6972 19320
rect 7104 19314 7156 19320
rect 7300 19334 7328 19654
rect 7300 19306 7420 19334
rect 7392 18902 7420 19306
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 17882 6960 18702
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6932 16114 6960 17818
rect 7024 17678 7052 18226
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7116 17542 7144 18022
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7208 17270 7236 18158
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17678 7420 17818
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 7208 16998 7236 17206
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 15706 6960 16050
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 12986 6960 13806
rect 7024 13394 7052 15302
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14278 7328 14894
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6380 12406 6776 12434
rect 6184 11892 6236 11898
rect 6012 11852 6184 11880
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5920 10130 5948 10678
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5814 9616 5870 9625
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5814 9551 5870 9560
rect 5724 9522 5776 9528
rect 5552 9110 5580 9522
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5540 8968 5592 8974
rect 5644 8956 5672 9522
rect 5736 9178 5764 9522
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5828 8974 5856 9551
rect 5592 8928 5672 8956
rect 5816 8968 5868 8974
rect 5540 8910 5592 8916
rect 5816 8910 5868 8916
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5828 7954 5856 8774
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7342 5856 7890
rect 5920 7886 5948 8774
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5460 6718 5580 6746
rect 5354 6695 5410 6704
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5368 6322 5396 6598
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5276 6174 5396 6202
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5778 5304 6054
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5368 3754 5396 6174
rect 5460 5642 5488 6598
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5552 5522 5580 6718
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5460 5494 5580 5522
rect 5460 4434 5488 5494
rect 5644 5114 5672 6258
rect 5736 6225 5764 6258
rect 5722 6216 5778 6225
rect 5722 6151 5778 6160
rect 5644 5086 5764 5114
rect 5736 5030 5764 5086
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4622 5764 4966
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5460 4406 5580 4434
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5276 3738 5396 3754
rect 5264 3732 5396 3738
rect 5316 3726 5396 3732
rect 5264 3674 5316 3680
rect 5460 2922 5488 4218
rect 5552 4146 5580 4406
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 6012 4078 6040 11852
rect 6184 11834 6236 11840
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6104 9586 6132 10474
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6104 8022 6132 9522
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7818 6132 7958
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 6934 6132 7346
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6196 6322 6224 10134
rect 6288 9722 6316 11562
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 6866 6316 8978
rect 6380 7206 6408 12406
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6564 11354 6592 11698
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10538 6592 11154
rect 6656 11150 6684 11494
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10742 6684 11086
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6748 10538 6776 11698
rect 6840 11354 6868 11698
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6932 10470 6960 11086
rect 7116 10606 7144 14010
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7208 13258 7236 13398
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 10742 7236 11290
rect 7300 11150 7328 14214
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7392 13530 7420 13942
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6840 10282 6868 10406
rect 6840 10254 6960 10282
rect 6932 9994 6960 10254
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6550 7783 6606 7792
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6840 6934 6868 7754
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5846 6776 6054
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5828 2990 5856 3402
rect 6012 3194 6040 3878
rect 6748 3398 6776 5782
rect 6840 5370 6868 6870
rect 6932 6798 6960 7890
rect 7024 7478 7052 9522
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7116 7546 7144 7686
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7024 6458 7052 7142
rect 7116 6798 7144 7482
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7208 6458 7236 7686
rect 7300 7546 7328 8366
rect 7392 8090 7420 8434
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7484 7954 7512 24670
rect 7668 23474 7696 24822
rect 8128 24750 8156 25366
rect 8220 24818 8248 25434
rect 8312 25362 8340 25774
rect 8668 25774 8720 25780
rect 8574 25735 8630 25744
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 8312 24818 8340 25298
rect 8588 25294 8616 25638
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8588 24886 8616 25094
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 7668 23446 7788 23474
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 7576 22574 7604 23122
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 7576 22234 7604 22510
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 7668 21622 7696 23054
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7576 20874 7604 21354
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7668 20058 7696 20402
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7668 19514 7696 19790
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7576 18766 7604 19314
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7668 18290 7696 18838
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7576 17882 7604 18226
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 17202 7696 17614
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12986 7604 13126
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7668 12918 7696 14962
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7760 12434 7788 23446
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7852 21010 7880 21490
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7852 20777 7880 20946
rect 7838 20768 7894 20777
rect 7838 20703 7894 20712
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 18834 7880 20402
rect 8036 18970 8064 22578
rect 8128 22094 8156 24686
rect 8680 24410 8708 25774
rect 8944 25696 8996 25702
rect 8944 25638 8996 25644
rect 8956 25294 8984 25638
rect 9048 25498 9076 25910
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8944 25288 8996 25294
rect 8944 25230 8996 25236
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8404 23730 8432 24142
rect 8758 23760 8814 23769
rect 8392 23724 8444 23730
rect 8758 23695 8814 23704
rect 8392 23666 8444 23672
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8220 22506 8248 22714
rect 8208 22500 8260 22506
rect 8208 22442 8260 22448
rect 8680 22166 8708 23462
rect 8668 22160 8720 22166
rect 8668 22102 8720 22108
rect 8128 22066 8248 22094
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7852 18737 7880 18770
rect 7838 18728 7894 18737
rect 7838 18663 7894 18672
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17746 7972 18022
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17134 7972 17478
rect 8036 17320 8064 18158
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8128 17882 8156 18022
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8036 17292 8156 17320
rect 8024 17196 8076 17202
rect 8128 17184 8156 17292
rect 8220 17252 8248 22066
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8312 20942 8340 21966
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 19514 8340 20878
rect 8404 20466 8432 21626
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8404 20058 8432 20198
rect 8482 20088 8538 20097
rect 8392 20052 8444 20058
rect 8482 20023 8538 20032
rect 8392 19994 8444 20000
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8496 19310 8524 20023
rect 8588 19446 8616 20742
rect 8680 20398 8708 22102
rect 8772 22030 8800 23695
rect 8864 23186 8892 24754
rect 9692 24721 9720 26182
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10152 25498 10180 25910
rect 10244 25906 10272 26250
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10230 25596 10538 25605
rect 10230 25594 10236 25596
rect 10292 25594 10316 25596
rect 10372 25594 10396 25596
rect 10452 25594 10476 25596
rect 10532 25594 10538 25596
rect 10292 25542 10294 25594
rect 10474 25542 10476 25594
rect 10230 25540 10236 25542
rect 10292 25540 10316 25542
rect 10372 25540 10396 25542
rect 10452 25540 10476 25542
rect 10532 25540 10538 25542
rect 10230 25531 10538 25540
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10414 25392 10470 25401
rect 10414 25327 10416 25336
rect 10468 25327 10470 25336
rect 10416 25298 10468 25304
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 10508 25220 10560 25226
rect 10612 25208 10640 25638
rect 10560 25180 10640 25208
rect 10508 25162 10560 25168
rect 9678 24712 9734 24721
rect 9678 24647 9734 24656
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 8864 22030 8892 23122
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22030 8984 22374
rect 9140 22030 9168 24142
rect 9692 23882 9720 24550
rect 9784 24138 9812 25162
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9646 23866 9720 23882
rect 9634 23860 9720 23866
rect 9686 23854 9720 23860
rect 9770 23896 9826 23905
rect 9770 23831 9772 23840
rect 9634 23802 9686 23808
rect 9824 23831 9826 23840
rect 10152 23848 10180 25094
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10230 24508 10538 24517
rect 10230 24506 10236 24508
rect 10292 24506 10316 24508
rect 10372 24506 10396 24508
rect 10452 24506 10476 24508
rect 10532 24506 10538 24508
rect 10292 24454 10294 24506
rect 10474 24454 10476 24506
rect 10230 24452 10236 24454
rect 10292 24452 10316 24454
rect 10372 24452 10396 24454
rect 10452 24452 10476 24454
rect 10532 24452 10538 24454
rect 10230 24443 10538 24452
rect 10612 24410 10640 24754
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10506 23896 10562 23905
rect 10152 23820 10456 23848
rect 10506 23831 10562 23840
rect 9772 23802 9824 23808
rect 10138 23760 10194 23769
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9772 23724 9824 23730
rect 10138 23695 10194 23704
rect 10324 23724 10376 23730
rect 9772 23666 9824 23672
rect 9508 23168 9536 23666
rect 9784 23526 9812 23666
rect 10152 23662 10180 23695
rect 10324 23666 10376 23672
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10048 23588 10100 23594
rect 10048 23530 10100 23536
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9784 23322 9812 23462
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9588 23180 9640 23186
rect 9508 23140 9588 23168
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 9232 22778 9260 22986
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8772 19854 8800 21966
rect 8864 21690 8892 21966
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8850 20360 8906 20369
rect 8850 20295 8906 20304
rect 8864 20262 8892 20295
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8956 20040 8984 20878
rect 9036 20052 9088 20058
rect 8956 20012 9036 20040
rect 9036 19994 9088 20000
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8760 19848 8812 19854
rect 9140 19802 9168 21966
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9218 20224 9274 20233
rect 9218 20159 9274 20168
rect 9232 20058 9260 20159
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9324 19854 9352 20334
rect 8760 19790 8812 19796
rect 8680 19666 8708 19790
rect 8864 19774 9168 19802
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 8864 19666 8892 19774
rect 8680 19638 8892 19666
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8392 19304 8444 19310
rect 8298 19272 8354 19281
rect 8392 19246 8444 19252
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8298 19207 8354 19216
rect 8312 18902 8340 19207
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17678 8340 18022
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8404 17542 8432 19246
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8392 17264 8444 17270
rect 8220 17224 8392 17252
rect 8392 17206 8444 17212
rect 8128 17156 8248 17184
rect 8024 17138 8076 17144
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8036 17082 8064 17138
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 16250 7880 16390
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 15638 7972 17070
rect 8036 17054 8156 17082
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16250 8064 16458
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8128 15450 8156 17054
rect 8220 16980 8248 17156
rect 8392 16992 8444 16998
rect 8220 16952 8392 16980
rect 8392 16934 8444 16940
rect 8208 15496 8260 15502
rect 8128 15444 8208 15450
rect 8128 15438 8260 15444
rect 8128 15422 8248 15438
rect 8220 14482 8248 15422
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 7852 12646 7880 14282
rect 8128 13802 8156 14282
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8128 13394 8156 13738
rect 8404 13734 8432 16934
rect 8496 16590 8524 18770
rect 8680 18290 8708 18838
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8588 17338 8616 17614
rect 8772 17338 8800 17614
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16590 8616 17002
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8760 16584 8812 16590
rect 8864 16572 8892 19638
rect 8956 18426 8984 19654
rect 9048 18834 9076 19654
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 9048 17882 9076 18634
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9048 17678 9076 17818
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8812 16544 8892 16572
rect 8944 16584 8996 16590
rect 8760 16526 8812 16532
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8496 14958 8524 15438
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8588 14278 8616 16186
rect 8864 15065 8892 16544
rect 8942 16552 8944 16561
rect 8996 16552 8998 16561
rect 8942 16487 8998 16496
rect 9140 15502 9168 19246
rect 9232 18426 9260 19790
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9324 16572 9352 19790
rect 9508 18970 9536 23140
rect 9588 23122 9640 23128
rect 9968 23050 9996 23462
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9770 22808 9826 22817
rect 9770 22743 9826 22752
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9600 21554 9628 21830
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9692 21486 9720 22510
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9692 20874 9720 21422
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 20602 9628 20742
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9692 18306 9720 19994
rect 9784 19174 9812 22743
rect 10060 22250 10088 23530
rect 10336 23508 10364 23666
rect 10428 23594 10456 23820
rect 10520 23662 10548 23831
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 10152 23480 10364 23508
rect 10152 22778 10180 23480
rect 10230 23420 10538 23429
rect 10230 23418 10236 23420
rect 10292 23418 10316 23420
rect 10372 23418 10396 23420
rect 10452 23418 10476 23420
rect 10532 23418 10538 23420
rect 10292 23366 10294 23418
rect 10474 23366 10476 23418
rect 10230 23364 10236 23366
rect 10292 23364 10316 23366
rect 10372 23364 10396 23366
rect 10452 23364 10476 23366
rect 10532 23364 10538 23366
rect 10230 23355 10538 23364
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10140 22500 10192 22506
rect 10140 22442 10192 22448
rect 9876 22222 10088 22250
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9232 16544 9352 16572
rect 9416 18278 9720 18306
rect 9232 16250 9260 16544
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9324 15706 9352 16050
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8850 15056 8906 15065
rect 8850 14991 8906 15000
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8312 13462 8340 13670
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8128 13297 8156 13330
rect 8404 13326 8432 13670
rect 8392 13320 8444 13326
rect 8114 13288 8170 13297
rect 8392 13262 8444 13268
rect 8114 13223 8170 13232
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12850 8156 13126
rect 8588 12986 8616 14214
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 13530 8800 13806
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7760 12406 8064 12434
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7576 11898 7604 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 9654 7604 11018
rect 7760 10470 7788 11698
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7668 8090 7696 9998
rect 7760 9586 7788 10406
rect 7852 10146 7880 12174
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7944 10266 7972 10542
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7852 10118 7972 10146
rect 7944 10062 7972 10118
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7852 9722 7880 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 8634 7880 9522
rect 7944 9382 7972 9862
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7562 7512 7890
rect 7748 7880 7800 7886
rect 7654 7848 7710 7857
rect 7748 7822 7800 7828
rect 7654 7783 7710 7792
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7392 7534 7512 7562
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7392 6322 7420 7534
rect 7668 7410 7696 7783
rect 7760 7478 7788 7822
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7852 7274 7880 8230
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7838 7168 7894 7177
rect 7760 6882 7788 7142
rect 7838 7103 7894 7112
rect 7852 7002 7880 7103
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7760 6854 7880 6882
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7024 5778 7052 6258
rect 7392 5914 7420 6258
rect 7484 5914 7512 6666
rect 7576 6610 7604 6734
rect 7576 6582 7696 6610
rect 7668 6118 7696 6582
rect 7760 6458 7788 6734
rect 7852 6662 7880 6854
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7944 6225 7972 9318
rect 7930 6216 7986 6225
rect 7930 6151 7986 6160
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7576 5914 7604 6054
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7392 5642 7420 5850
rect 7668 5846 7696 6054
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 4826 7696 5170
rect 7944 4826 7972 5306
rect 8036 5030 8064 12406
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5816 2984 5868 2990
rect 6748 2972 6776 3334
rect 6840 3194 6868 3878
rect 7024 3738 7052 3878
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 3194 7144 3402
rect 7300 3194 7328 3878
rect 7392 3738 7420 4082
rect 7576 4078 7604 4422
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7852 3670 7880 4082
rect 7944 4010 7972 4150
rect 8036 4146 8064 4558
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7760 3058 7788 3470
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 6828 2984 6880 2990
rect 6748 2944 6828 2972
rect 5816 2926 5868 2932
rect 6828 2926 6880 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6564 2650 6592 2858
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 4068 2440 4120 2446
rect 3882 2408 3938 2417
rect 3882 2343 3884 2352
rect 3936 2343 3938 2352
rect 3988 2400 4068 2428
rect 3884 2314 3936 2320
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 1170 3464 2246
rect 3988 1306 4016 2400
rect 4068 2382 4120 2388
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 3252 1142 3464 1170
rect 3896 1278 4016 1306
rect 3252 800 3280 1142
rect 3896 800 3924 1278
rect 4632 1170 4660 2246
rect 4703 2204 5011 2213
rect 4703 2202 4709 2204
rect 4765 2202 4789 2204
rect 4845 2202 4869 2204
rect 4925 2202 4949 2204
rect 5005 2202 5011 2204
rect 4765 2150 4767 2202
rect 4947 2150 4949 2202
rect 4703 2148 4709 2150
rect 4765 2148 4789 2150
rect 4845 2148 4869 2150
rect 4925 2148 4949 2150
rect 5005 2148 5011 2150
rect 4703 2139 5011 2148
rect 5184 2106 5212 2314
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5276 1170 5304 2246
rect 5368 2038 5396 2314
rect 5460 2038 5488 2450
rect 6460 2440 6512 2446
rect 7196 2440 7248 2446
rect 6460 2382 6512 2388
rect 7116 2400 7196 2428
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 4540 1142 4660 1170
rect 5184 1142 5304 1170
rect 4540 800 4568 1142
rect 5184 800 5212 1142
rect 6472 800 6500 2382
rect 7116 800 7144 2400
rect 7840 2440 7892 2446
rect 7196 2382 7248 2388
rect 7760 2400 7840 2428
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 2106 7420 2246
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7760 800 7788 2400
rect 7840 2382 7892 2388
rect 8128 1970 8156 12786
rect 8220 11762 8248 12786
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8312 11694 8340 12854
rect 8588 12306 8616 12922
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11286 8340 11630
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 8906 8248 9998
rect 8312 9178 8340 11222
rect 8680 11150 8708 12922
rect 8864 11898 8892 14991
rect 9416 12646 9444 18278
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9508 17610 9536 18158
rect 9678 17776 9734 17785
rect 9678 17711 9680 17720
rect 9732 17711 9734 17720
rect 9680 17682 9732 17688
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9508 16250 9536 17546
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16658 9628 17002
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9600 13682 9628 15642
rect 9692 13818 9720 17546
rect 9784 14362 9812 18906
rect 9876 14532 9904 22222
rect 9954 22128 10010 22137
rect 10152 22098 10180 22442
rect 10230 22332 10538 22341
rect 10230 22330 10236 22332
rect 10292 22330 10316 22332
rect 10372 22330 10396 22332
rect 10452 22330 10476 22332
rect 10532 22330 10538 22332
rect 10292 22278 10294 22330
rect 10474 22278 10476 22330
rect 10230 22276 10236 22278
rect 10292 22276 10316 22278
rect 10372 22276 10396 22278
rect 10452 22276 10476 22278
rect 10532 22276 10538 22278
rect 10230 22267 10538 22276
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10244 22137 10272 22170
rect 10230 22128 10286 22137
rect 9954 22063 10010 22072
rect 10140 22092 10192 22098
rect 9968 21622 9996 22063
rect 10230 22063 10286 22072
rect 10140 22034 10192 22040
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 10046 21584 10102 21593
rect 10046 21519 10102 21528
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9968 20330 9996 20470
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9968 15706 9996 19110
rect 10060 17252 10088 21519
rect 10152 21350 10180 22034
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 21078 10180 21286
rect 10230 21244 10538 21253
rect 10230 21242 10236 21244
rect 10292 21242 10316 21244
rect 10372 21242 10396 21244
rect 10452 21242 10476 21244
rect 10532 21242 10538 21244
rect 10292 21190 10294 21242
rect 10474 21190 10476 21242
rect 10230 21188 10236 21190
rect 10292 21188 10316 21190
rect 10372 21188 10396 21190
rect 10452 21188 10476 21190
rect 10532 21188 10538 21190
rect 10230 21179 10538 21188
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10336 20806 10364 20878
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10152 20602 10180 20742
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 20058 10180 20198
rect 10230 20156 10538 20165
rect 10230 20154 10236 20156
rect 10292 20154 10316 20156
rect 10372 20154 10396 20156
rect 10452 20154 10476 20156
rect 10532 20154 10538 20156
rect 10292 20102 10294 20154
rect 10474 20102 10476 20154
rect 10230 20100 10236 20102
rect 10292 20100 10316 20102
rect 10372 20100 10396 20102
rect 10452 20100 10476 20102
rect 10532 20100 10538 20102
rect 10230 20091 10538 20100
rect 10704 20097 10732 26454
rect 12268 26382 12296 28381
rect 12912 26382 12940 28381
rect 14476 26586 14504 28478
rect 14830 28381 14886 29181
rect 15474 28381 15530 29181
rect 16762 28381 16818 29181
rect 17406 28381 17462 29181
rect 18050 28381 18106 29181
rect 18694 28506 18750 29181
rect 18694 28478 19104 28506
rect 18694 28381 18750 28478
rect 14464 26580 14516 26586
rect 14464 26522 14516 26528
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 14096 26308 14148 26314
rect 14096 26250 14148 26256
rect 10890 26140 11198 26149
rect 10890 26138 10896 26140
rect 10952 26138 10976 26140
rect 11032 26138 11056 26140
rect 11112 26138 11136 26140
rect 11192 26138 11198 26140
rect 10952 26086 10954 26138
rect 11134 26086 11136 26138
rect 10890 26084 10896 26086
rect 10952 26084 10976 26086
rect 11032 26084 11056 26086
rect 11112 26084 11136 26086
rect 11192 26084 11198 26086
rect 10890 26075 11198 26084
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10888 25140 10916 25774
rect 11428 25764 11480 25770
rect 11428 25706 11480 25712
rect 11440 25498 11468 25706
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 10796 25112 10916 25140
rect 11244 25152 11296 25158
rect 10796 24886 10824 25112
rect 11244 25094 11296 25100
rect 10890 25052 11198 25061
rect 10890 25050 10896 25052
rect 10952 25050 10976 25052
rect 11032 25050 11056 25052
rect 11112 25050 11136 25052
rect 11192 25050 11198 25052
rect 10952 24998 10954 25050
rect 11134 24998 11136 25050
rect 10890 24996 10896 24998
rect 10952 24996 10976 24998
rect 11032 24996 11056 24998
rect 11112 24996 11136 24998
rect 11192 24996 11198 24998
rect 10890 24987 11198 24996
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10876 24744 10928 24750
rect 10796 24704 10876 24732
rect 10796 22030 10824 24704
rect 10876 24686 10928 24692
rect 11256 24274 11284 25094
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10890 23964 11198 23973
rect 10890 23962 10896 23964
rect 10952 23962 10976 23964
rect 11032 23962 11056 23964
rect 11112 23962 11136 23964
rect 11192 23962 11198 23964
rect 10952 23910 10954 23962
rect 11134 23910 11136 23962
rect 10890 23908 10896 23910
rect 10952 23908 10976 23910
rect 11032 23908 11056 23910
rect 11112 23908 11136 23910
rect 11192 23908 11198 23910
rect 10890 23899 11198 23908
rect 10890 22876 11198 22885
rect 10890 22874 10896 22876
rect 10952 22874 10976 22876
rect 11032 22874 11056 22876
rect 11112 22874 11136 22876
rect 11192 22874 11198 22876
rect 10952 22822 10954 22874
rect 11134 22822 11136 22874
rect 10890 22820 10896 22822
rect 10952 22820 10976 22822
rect 11032 22820 11056 22822
rect 11112 22820 11136 22822
rect 11192 22820 11198 22822
rect 10890 22811 11198 22820
rect 11256 22642 11284 24210
rect 11348 24138 11376 24550
rect 11440 24410 11468 25434
rect 11532 25362 11560 25638
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 11808 25226 11836 25638
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11992 24954 12020 25842
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11532 24070 11560 24550
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11992 23798 12020 24754
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11348 22778 11376 22986
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 10784 22024 10836 22030
rect 10782 21992 10784 22001
rect 11336 22024 11388 22030
rect 10836 21992 10838 22001
rect 11336 21966 11388 21972
rect 10782 21927 10838 21936
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21622 10824 21830
rect 10890 21788 11198 21797
rect 10890 21786 10896 21788
rect 10952 21786 10976 21788
rect 11032 21786 11056 21788
rect 11112 21786 11136 21788
rect 11192 21786 11198 21788
rect 10952 21734 10954 21786
rect 11134 21734 11136 21786
rect 10890 21732 10896 21734
rect 10952 21732 10976 21734
rect 11032 21732 11056 21734
rect 11112 21732 11136 21734
rect 11192 21732 11198 21734
rect 10890 21723 11198 21732
rect 11348 21690 11376 21966
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10690 20088 10746 20097
rect 10140 20052 10192 20058
rect 10690 20023 10746 20032
rect 10140 19994 10192 20000
rect 10704 19514 10732 20023
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10230 19068 10538 19077
rect 10230 19066 10236 19068
rect 10292 19066 10316 19068
rect 10372 19066 10396 19068
rect 10452 19066 10476 19068
rect 10532 19066 10538 19068
rect 10292 19014 10294 19066
rect 10474 19014 10476 19066
rect 10230 19012 10236 19014
rect 10292 19012 10316 19014
rect 10372 19012 10396 19014
rect 10452 19012 10476 19014
rect 10532 19012 10538 19014
rect 10230 19003 10538 19012
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10152 18426 10180 18634
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10230 17980 10538 17989
rect 10230 17978 10236 17980
rect 10292 17978 10316 17980
rect 10372 17978 10396 17980
rect 10452 17978 10476 17980
rect 10532 17978 10538 17980
rect 10292 17926 10294 17978
rect 10474 17926 10476 17978
rect 10230 17924 10236 17926
rect 10292 17924 10316 17926
rect 10372 17924 10396 17926
rect 10452 17924 10476 17926
rect 10532 17924 10538 17926
rect 10230 17915 10538 17924
rect 10612 17882 10640 18634
rect 10704 18426 10732 19110
rect 10796 18850 10824 21558
rect 11440 21146 11468 21898
rect 11624 21146 11652 22034
rect 11808 22030 11836 23734
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11440 20942 11468 21082
rect 11796 21072 11848 21078
rect 11716 21032 11796 21060
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 10890 20700 11198 20709
rect 10890 20698 10896 20700
rect 10952 20698 10976 20700
rect 11032 20698 11056 20700
rect 11112 20698 11136 20700
rect 11192 20698 11198 20700
rect 10952 20646 10954 20698
rect 11134 20646 11136 20698
rect 10890 20644 10896 20646
rect 10952 20644 10976 20646
rect 11032 20644 11056 20646
rect 11112 20644 11136 20646
rect 11192 20644 11198 20646
rect 10890 20635 11198 20644
rect 11152 20460 11204 20466
rect 11256 20448 11284 20810
rect 11532 20466 11560 20810
rect 11204 20420 11284 20448
rect 11520 20460 11572 20466
rect 11152 20402 11204 20408
rect 11520 20402 11572 20408
rect 11164 20058 11192 20402
rect 11716 20369 11744 21032
rect 11796 21014 11848 21020
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 20602 11928 20810
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11702 20360 11758 20369
rect 11428 20324 11480 20330
rect 11702 20295 11758 20304
rect 11428 20266 11480 20272
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11348 19990 11376 20198
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11440 19854 11468 20266
rect 11716 20262 11744 20295
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 10890 19612 11198 19621
rect 10890 19610 10896 19612
rect 10952 19610 10976 19612
rect 11032 19610 11056 19612
rect 11112 19610 11136 19612
rect 11192 19610 11198 19612
rect 10952 19558 10954 19610
rect 11134 19558 11136 19610
rect 10890 19556 10896 19558
rect 10952 19556 10976 19558
rect 11032 19556 11056 19558
rect 11112 19556 11136 19558
rect 11192 19556 11198 19558
rect 10890 19547 11198 19556
rect 10966 18864 11022 18873
rect 10796 18822 10966 18850
rect 11348 18834 11376 19790
rect 10966 18799 11022 18808
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 10890 18524 11198 18533
rect 10890 18522 10896 18524
rect 10952 18522 10976 18524
rect 11032 18522 11056 18524
rect 11112 18522 11136 18524
rect 11192 18522 11198 18524
rect 10952 18470 10954 18522
rect 11134 18470 11136 18522
rect 10890 18468 10896 18470
rect 10952 18468 10976 18470
rect 11032 18468 11056 18470
rect 11112 18468 11136 18470
rect 11192 18468 11198 18470
rect 10890 18459 11198 18468
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 11348 18222 11376 18770
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10060 17224 10180 17252
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 15910 10088 16390
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 15162 9996 15438
rect 10060 15366 10088 15846
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10048 14544 10100 14550
rect 9876 14504 9996 14532
rect 9784 14334 9904 14362
rect 9772 13864 9824 13870
rect 9692 13812 9772 13818
rect 9692 13806 9824 13812
rect 9692 13790 9812 13806
rect 9600 13654 9720 13682
rect 9692 13274 9720 13654
rect 9784 13394 9812 13790
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9770 13288 9826 13297
rect 9692 13246 9770 13274
rect 9770 13223 9826 13232
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12850 9812 13126
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9680 12776 9732 12782
rect 9876 12730 9904 14334
rect 9680 12718 9732 12724
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 9416 11676 9444 12242
rect 9508 11778 9536 12650
rect 9692 12238 9720 12718
rect 9784 12702 9904 12730
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11898 9628 12038
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9680 11824 9732 11830
rect 9508 11772 9680 11778
rect 9508 11766 9732 11772
rect 9508 11750 9720 11766
rect 9416 11648 9628 11676
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11354 9444 11494
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10062 8432 10950
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10266 8524 10678
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8404 8498 8432 9522
rect 8588 9110 8616 9522
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 9042 8708 11086
rect 8772 10810 8800 11086
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8772 9586 8800 10746
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9654 9352 9862
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9324 8634 9352 8910
rect 9416 8838 9444 9998
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8220 7750 8248 7958
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 7177 8248 7346
rect 8312 7274 8340 7890
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7268 8352 7274
rect 8404 7256 8432 7482
rect 8496 7324 8524 7822
rect 8680 7546 8708 7958
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8588 7426 8616 7482
rect 8588 7398 8708 7426
rect 8680 7342 8708 7398
rect 8772 7342 8800 8026
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8576 7336 8628 7342
rect 8496 7296 8576 7324
rect 8576 7278 8628 7284
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8404 7228 8524 7256
rect 8300 7210 8352 7216
rect 8206 7168 8262 7177
rect 8206 7103 8262 7112
rect 8496 6984 8524 7228
rect 8404 6956 8524 6984
rect 8404 6798 8432 6956
rect 8588 6882 8616 7278
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 7002 8708 7142
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8496 6854 8616 6882
rect 8772 6866 8800 7278
rect 8864 7002 8892 7822
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7546 8984 7686
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9140 7426 9168 7822
rect 9048 7410 9168 7426
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9036 7404 9168 7410
rect 9088 7398 9168 7404
rect 9036 7346 9088 7352
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8760 6860 8812 6866
rect 8496 6798 8524 6854
rect 8760 6802 8812 6808
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6458 8340 6666
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 6390 8432 6734
rect 8772 6458 8800 6802
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8404 5370 8432 6326
rect 8772 5914 8800 6394
rect 8864 6338 8892 6938
rect 9048 6730 9076 7346
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 7002 9168 7142
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9140 6458 9168 6734
rect 9232 6458 9260 6938
rect 9324 6798 9352 7414
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9416 6730 9444 6870
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8864 6322 8984 6338
rect 8864 6316 8996 6322
rect 8864 6310 8944 6316
rect 8944 6258 8996 6264
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 5574 8984 6258
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4078 9076 4966
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8220 3738 8248 4014
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3602 8340 4014
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3602 8432 3878
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8312 3194 8340 3538
rect 8956 3194 8984 3946
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9140 2650 9168 3402
rect 9416 3398 9444 5782
rect 9508 5302 9536 10610
rect 9600 9110 9628 11648
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9692 9217 9720 10746
rect 9784 9489 9812 12702
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9678 9208 9734 9217
rect 9784 9178 9812 9318
rect 9678 9143 9734 9152
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9588 9104 9640 9110
rect 9876 9081 9904 12582
rect 9588 9046 9640 9052
rect 9862 9072 9918 9081
rect 9968 9058 9996 14504
rect 10048 14486 10100 14492
rect 10060 14006 10088 14486
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10060 12306 10088 13330
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11354 10088 12038
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10152 10810 10180 17224
rect 10230 16892 10538 16901
rect 10230 16890 10236 16892
rect 10292 16890 10316 16892
rect 10372 16890 10396 16892
rect 10452 16890 10476 16892
rect 10532 16890 10538 16892
rect 10292 16838 10294 16890
rect 10474 16838 10476 16890
rect 10230 16836 10236 16838
rect 10292 16836 10316 16838
rect 10372 16836 10396 16838
rect 10452 16836 10476 16838
rect 10532 16836 10538 16838
rect 10230 16827 10538 16836
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 16046 10456 16594
rect 10506 16552 10562 16561
rect 10506 16487 10562 16496
rect 10520 16114 10548 16487
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10612 15978 10640 16662
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 16028 10732 16458
rect 10796 16250 10824 17614
rect 10890 17436 11198 17445
rect 10890 17434 10896 17436
rect 10952 17434 10976 17436
rect 11032 17434 11056 17436
rect 11112 17434 11136 17436
rect 11192 17434 11198 17436
rect 10952 17382 10954 17434
rect 11134 17382 11136 17434
rect 10890 17380 10896 17382
rect 10952 17380 10976 17382
rect 11032 17380 11056 17382
rect 11112 17380 11136 17382
rect 11192 17380 11198 17382
rect 10890 17371 11198 17380
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 16794 11100 17138
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16794 11192 16934
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11348 16522 11376 18158
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 10890 16348 11198 16357
rect 10890 16346 10896 16348
rect 10952 16346 10976 16348
rect 11032 16346 11056 16348
rect 11112 16346 11136 16348
rect 11192 16346 11198 16348
rect 10952 16294 10954 16346
rect 11134 16294 11136 16346
rect 10890 16292 10896 16294
rect 10952 16292 10976 16294
rect 11032 16292 11056 16294
rect 11112 16292 11136 16294
rect 11192 16292 11198 16294
rect 10890 16283 11198 16292
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10876 16040 10928 16046
rect 10704 16000 10876 16028
rect 10876 15982 10928 15988
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10230 15804 10538 15813
rect 10230 15802 10236 15804
rect 10292 15802 10316 15804
rect 10372 15802 10396 15804
rect 10452 15802 10476 15804
rect 10532 15802 10538 15804
rect 10292 15750 10294 15802
rect 10474 15750 10476 15802
rect 10230 15748 10236 15750
rect 10292 15748 10316 15750
rect 10372 15748 10396 15750
rect 10452 15748 10476 15750
rect 10532 15748 10538 15750
rect 10230 15739 10538 15748
rect 10230 14716 10538 14725
rect 10230 14714 10236 14716
rect 10292 14714 10316 14716
rect 10372 14714 10396 14716
rect 10452 14714 10476 14716
rect 10532 14714 10538 14716
rect 10292 14662 10294 14714
rect 10474 14662 10476 14714
rect 10230 14660 10236 14662
rect 10292 14660 10316 14662
rect 10372 14660 10396 14662
rect 10452 14660 10476 14662
rect 10532 14660 10538 14662
rect 10230 14651 10538 14660
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 14074 10364 14282
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10520 14006 10548 14350
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10520 13841 10548 13942
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10230 13628 10538 13637
rect 10230 13626 10236 13628
rect 10292 13626 10316 13628
rect 10372 13626 10396 13628
rect 10452 13626 10476 13628
rect 10532 13626 10538 13628
rect 10292 13574 10294 13626
rect 10474 13574 10476 13626
rect 10230 13572 10236 13574
rect 10292 13572 10316 13574
rect 10372 13572 10396 13574
rect 10452 13572 10476 13574
rect 10532 13572 10538 13574
rect 10230 13563 10538 13572
rect 10612 13530 10640 15914
rect 10888 15706 10916 15982
rect 10876 15700 10928 15706
rect 10796 15660 10876 15688
rect 10796 14958 10824 15660
rect 10876 15642 10928 15648
rect 10980 15502 11008 16186
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15502 11100 16050
rect 11348 16046 11376 16458
rect 11426 16416 11482 16425
rect 11426 16351 11482 16360
rect 11440 16182 11468 16351
rect 11532 16182 11560 19994
rect 11900 19922 11928 20402
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11624 18970 11652 19178
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11992 18766 12020 19110
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11808 18222 11836 18566
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11886 17640 11942 17649
rect 11704 17604 11756 17610
rect 11886 17575 11942 17584
rect 11704 17546 11756 17552
rect 11716 16250 11744 17546
rect 11900 17270 11928 17575
rect 11888 17264 11940 17270
rect 11808 17224 11888 17252
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11520 16176 11572 16182
rect 11572 16136 11652 16164
rect 11520 16118 11572 16124
rect 11336 16040 11388 16046
rect 11242 16008 11298 16017
rect 11152 15972 11204 15978
rect 11336 15982 11388 15988
rect 11242 15943 11298 15952
rect 11152 15914 11204 15920
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11164 15366 11192 15914
rect 11256 15570 11284 15943
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 15570 11376 15846
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11624 15502 11652 16136
rect 11808 16114 11836 17224
rect 11888 17206 11940 17212
rect 11992 17116 12020 18566
rect 12084 17898 12112 26250
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12176 24410 12204 24618
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12176 24313 12204 24346
rect 12162 24304 12218 24313
rect 12162 24239 12218 24248
rect 12268 24138 12296 24550
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12452 23866 12480 24754
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12256 23588 12308 23594
rect 12256 23530 12308 23536
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12176 22778 12204 22918
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12268 22234 12296 23530
rect 12636 23202 12664 26182
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12808 25424 12860 25430
rect 12808 25366 12860 25372
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12728 24886 12756 25162
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12820 24682 12848 25366
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12820 23594 12848 24618
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12912 23474 12940 25434
rect 13188 25378 13216 26182
rect 12820 23446 12940 23474
rect 13004 25350 13216 25378
rect 13820 25424 13872 25430
rect 13820 25366 13872 25372
rect 13728 25356 13780 25362
rect 12636 23174 12756 23202
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12636 22778 12664 23054
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 12360 22234 12388 22646
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12164 22094 12216 22098
rect 12268 22094 12296 22170
rect 12164 22092 12296 22094
rect 12216 22066 12296 22092
rect 12164 22034 12216 22040
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12268 20330 12296 21490
rect 12360 20590 12572 20618
rect 12728 20602 12756 23174
rect 12820 21486 12848 23446
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12360 19310 12388 20590
rect 12544 20516 12572 20590
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12544 20488 12664 20516
rect 12636 20398 12664 20488
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 20058 12480 20198
rect 12544 20058 12572 20334
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12348 19304 12400 19310
rect 12346 19272 12348 19281
rect 12400 19272 12402 19281
rect 12346 19207 12402 19216
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12084 17870 12296 17898
rect 12072 17128 12124 17134
rect 11992 17088 12072 17116
rect 12072 17070 12124 17076
rect 12084 16658 12112 17070
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11612 15496 11664 15502
rect 11440 15456 11612 15484
rect 11152 15360 11204 15366
rect 11204 15320 11284 15348
rect 11152 15302 11204 15308
rect 10890 15260 11198 15269
rect 10890 15258 10896 15260
rect 10952 15258 10976 15260
rect 11032 15258 11056 15260
rect 11112 15258 11136 15260
rect 11192 15258 11198 15260
rect 10952 15206 10954 15258
rect 11134 15206 11136 15258
rect 10890 15204 10896 15206
rect 10952 15204 10976 15206
rect 11032 15204 11056 15206
rect 11112 15204 11136 15206
rect 11192 15204 11198 15206
rect 10890 15195 11198 15204
rect 11256 15144 11284 15320
rect 11072 15116 11284 15144
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 11072 14890 11100 15116
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10704 13802 10732 14826
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10796 13938 10824 14282
rect 10890 14172 11198 14181
rect 10890 14170 10896 14172
rect 10952 14170 10976 14172
rect 11032 14170 11056 14172
rect 11112 14170 11136 14172
rect 11192 14170 11198 14172
rect 10952 14118 10954 14170
rect 11134 14118 11136 14170
rect 10890 14116 10896 14118
rect 10952 14116 10976 14118
rect 11032 14116 11056 14118
rect 11112 14116 11136 14118
rect 11192 14116 11198 14118
rect 10890 14107 11198 14116
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 11256 13870 11284 14758
rect 11244 13864 11296 13870
rect 10782 13832 10838 13841
rect 10692 13796 10744 13802
rect 11244 13806 11296 13812
rect 10782 13767 10838 13776
rect 10692 13738 10744 13744
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10796 13326 10824 13767
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 12850 10732 13194
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10508 12776 10560 12782
rect 10560 12724 10640 12730
rect 10508 12718 10640 12724
rect 10520 12702 10640 12718
rect 10230 12540 10538 12549
rect 10230 12538 10236 12540
rect 10292 12538 10316 12540
rect 10372 12538 10396 12540
rect 10452 12538 10476 12540
rect 10532 12538 10538 12540
rect 10292 12486 10294 12538
rect 10474 12486 10476 12538
rect 10230 12484 10236 12486
rect 10292 12484 10316 12486
rect 10372 12484 10396 12486
rect 10452 12484 10476 12486
rect 10532 12484 10538 12486
rect 10230 12475 10538 12484
rect 10230 11452 10538 11461
rect 10230 11450 10236 11452
rect 10292 11450 10316 11452
rect 10372 11450 10396 11452
rect 10452 11450 10476 11452
rect 10532 11450 10538 11452
rect 10292 11398 10294 11450
rect 10474 11398 10476 11450
rect 10230 11396 10236 11398
rect 10292 11396 10316 11398
rect 10372 11396 10396 11398
rect 10452 11396 10476 11398
rect 10532 11396 10538 11398
rect 10230 11387 10538 11396
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10230 10364 10538 10373
rect 10230 10362 10236 10364
rect 10292 10362 10316 10364
rect 10372 10362 10396 10364
rect 10452 10362 10476 10364
rect 10532 10362 10538 10364
rect 10292 10310 10294 10362
rect 10474 10310 10476 10362
rect 10230 10308 10236 10310
rect 10292 10308 10316 10310
rect 10372 10308 10396 10310
rect 10452 10308 10476 10310
rect 10532 10308 10538 10310
rect 10230 10299 10538 10308
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9450 10180 9998
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 9654 10456 9862
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10230 9276 10538 9285
rect 10230 9274 10236 9276
rect 10292 9274 10316 9276
rect 10372 9274 10396 9276
rect 10452 9274 10476 9276
rect 10532 9274 10538 9276
rect 10292 9222 10294 9274
rect 10474 9222 10476 9274
rect 10230 9220 10236 9222
rect 10292 9220 10316 9222
rect 10372 9220 10396 9222
rect 10452 9220 10476 9222
rect 10532 9220 10538 9222
rect 10230 9211 10538 9220
rect 10138 9072 10194 9081
rect 9968 9030 10088 9058
rect 9862 9007 9918 9016
rect 9678 8936 9734 8945
rect 9678 8871 9734 8880
rect 9692 8566 9720 8871
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9600 6769 9628 8434
rect 9692 7562 9720 8502
rect 9784 8090 9812 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9692 7534 9812 7562
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9586 6760 9642 6769
rect 9586 6695 9642 6704
rect 9600 6322 9628 6695
rect 9692 6662 9720 7414
rect 9784 6798 9812 7534
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9678 6352 9734 6361
rect 9588 6316 9640 6322
rect 9876 6322 9904 7142
rect 9678 6287 9680 6296
rect 9588 6258 9640 6264
rect 9732 6287 9734 6296
rect 9864 6316 9916 6322
rect 9680 6258 9732 6264
rect 9864 6258 9916 6264
rect 9586 6216 9642 6225
rect 9642 6186 9720 6202
rect 9642 6180 9732 6186
rect 9642 6174 9680 6180
rect 9586 6151 9642 6160
rect 9680 6122 9732 6128
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4434 9812 4558
rect 9600 4406 9812 4434
rect 9600 4214 9628 4406
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3466 9904 3878
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9324 2990 9352 3334
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9416 2854 9444 3334
rect 9600 3058 9628 3402
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 3126 9812 3334
rect 10060 3194 10088 9030
rect 10138 9007 10194 9016
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9772 2984 9824 2990
rect 9862 2952 9918 2961
rect 9824 2932 9862 2938
rect 9772 2926 9862 2932
rect 9784 2910 9862 2926
rect 9862 2887 9918 2896
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 10152 2446 10180 9007
rect 10230 8188 10538 8197
rect 10230 8186 10236 8188
rect 10292 8186 10316 8188
rect 10372 8186 10396 8188
rect 10452 8186 10476 8188
rect 10532 8186 10538 8188
rect 10292 8134 10294 8186
rect 10474 8134 10476 8186
rect 10230 8132 10236 8134
rect 10292 8132 10316 8134
rect 10372 8132 10396 8134
rect 10452 8132 10476 8134
rect 10532 8132 10538 8134
rect 10230 8123 10538 8132
rect 10230 7100 10538 7109
rect 10230 7098 10236 7100
rect 10292 7098 10316 7100
rect 10372 7098 10396 7100
rect 10452 7098 10476 7100
rect 10532 7098 10538 7100
rect 10292 7046 10294 7098
rect 10474 7046 10476 7098
rect 10230 7044 10236 7046
rect 10292 7044 10316 7046
rect 10372 7044 10396 7046
rect 10452 7044 10476 7046
rect 10532 7044 10538 7046
rect 10230 7035 10538 7044
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 6118 10272 6258
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10230 6012 10538 6021
rect 10230 6010 10236 6012
rect 10292 6010 10316 6012
rect 10372 6010 10396 6012
rect 10452 6010 10476 6012
rect 10532 6010 10538 6012
rect 10292 5958 10294 6010
rect 10474 5958 10476 6010
rect 10230 5956 10236 5958
rect 10292 5956 10316 5958
rect 10372 5956 10396 5958
rect 10452 5956 10476 5958
rect 10532 5956 10538 5958
rect 10230 5947 10538 5956
rect 10230 4924 10538 4933
rect 10230 4922 10236 4924
rect 10292 4922 10316 4924
rect 10372 4922 10396 4924
rect 10452 4922 10476 4924
rect 10532 4922 10538 4924
rect 10292 4870 10294 4922
rect 10474 4870 10476 4922
rect 10230 4868 10236 4870
rect 10292 4868 10316 4870
rect 10372 4868 10396 4870
rect 10452 4868 10476 4870
rect 10532 4868 10538 4870
rect 10230 4859 10538 4868
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4214 10364 4422
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10230 3836 10538 3845
rect 10230 3834 10236 3836
rect 10292 3834 10316 3836
rect 10372 3834 10396 3836
rect 10452 3834 10476 3836
rect 10532 3834 10538 3836
rect 10292 3782 10294 3834
rect 10474 3782 10476 3834
rect 10230 3780 10236 3782
rect 10292 3780 10316 3782
rect 10372 3780 10396 3782
rect 10452 3780 10476 3782
rect 10532 3780 10538 3782
rect 10230 3771 10538 3780
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10520 3126 10548 3470
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10230 2748 10538 2757
rect 10230 2746 10236 2748
rect 10292 2746 10316 2748
rect 10372 2746 10396 2748
rect 10452 2746 10476 2748
rect 10532 2746 10538 2748
rect 10292 2694 10294 2746
rect 10474 2694 10476 2746
rect 10230 2692 10236 2694
rect 10292 2692 10316 2694
rect 10372 2692 10396 2694
rect 10452 2692 10476 2694
rect 10532 2692 10538 2694
rect 10230 2683 10538 2692
rect 10612 2650 10640 12702
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10704 11558 10732 12242
rect 10796 12238 10824 13262
rect 10890 13084 11198 13093
rect 10890 13082 10896 13084
rect 10952 13082 10976 13084
rect 11032 13082 11056 13084
rect 11112 13082 11136 13084
rect 11192 13082 11198 13084
rect 10952 13030 10954 13082
rect 11134 13030 11136 13082
rect 10890 13028 10896 13030
rect 10952 13028 10976 13030
rect 11032 13028 11056 13030
rect 11112 13028 11136 13030
rect 11192 13028 11198 13030
rect 10890 13019 11198 13028
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10980 12646 11008 12922
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11256 12646 11284 12854
rect 11440 12850 11468 15456
rect 11612 15438 11664 15444
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14346 11560 14758
rect 11900 14618 11928 16118
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13938 11652 14214
rect 11900 14074 11928 14554
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11704 13864 11756 13870
rect 11518 13832 11574 13841
rect 11704 13806 11756 13812
rect 11518 13767 11574 13776
rect 11612 13796 11664 13802
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10888 12374 10916 12582
rect 11532 12442 11560 13767
rect 11612 13738 11664 13744
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 11058 12336 11114 12345
rect 11624 12322 11652 13738
rect 11058 12271 11114 12280
rect 11256 12294 11652 12322
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10796 10810 10824 12174
rect 11072 12170 11100 12271
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10890 11996 11198 12005
rect 10890 11994 10896 11996
rect 10952 11994 10976 11996
rect 11032 11994 11056 11996
rect 11112 11994 11136 11996
rect 11192 11994 11198 11996
rect 10952 11942 10954 11994
rect 11134 11942 11136 11994
rect 10890 11940 10896 11942
rect 10952 11940 10976 11942
rect 11032 11940 11056 11942
rect 11112 11940 11136 11942
rect 11192 11940 11198 11942
rect 10890 11931 11198 11940
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 11014 11100 11086
rect 11164 11014 11192 11698
rect 11256 11642 11284 12294
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11898 11376 12038
rect 11716 11898 11744 13806
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11532 11762 11560 11834
rect 11520 11756 11572 11762
rect 11440 11716 11520 11744
rect 11256 11614 11376 11642
rect 11348 11218 11376 11614
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10890 10908 11198 10917
rect 10890 10906 10896 10908
rect 10952 10906 10976 10908
rect 11032 10906 11056 10908
rect 11112 10906 11136 10908
rect 11192 10906 11198 10908
rect 10952 10854 10954 10906
rect 11134 10854 11136 10906
rect 10890 10852 10896 10854
rect 10952 10852 10976 10854
rect 11032 10852 11056 10854
rect 11112 10852 11136 10854
rect 11192 10852 11198 10854
rect 10890 10843 11198 10852
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11256 10266 11284 11086
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11348 10198 11376 11154
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 10890 9820 11198 9829
rect 10890 9818 10896 9820
rect 10952 9818 10976 9820
rect 11032 9818 11056 9820
rect 11112 9818 11136 9820
rect 11192 9818 11198 9820
rect 10952 9766 10954 9818
rect 11134 9766 11136 9818
rect 10890 9764 10896 9766
rect 10952 9764 10976 9766
rect 11032 9764 11056 9766
rect 11112 9764 11136 9766
rect 11192 9764 11198 9766
rect 10890 9755 11198 9764
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 11152 9580 11204 9586
rect 11072 9518 11100 9551
rect 11152 9522 11204 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10782 9344 10838 9353
rect 10704 6322 10732 9318
rect 10782 9279 10838 9288
rect 10796 8566 10824 9279
rect 11164 9042 11192 9522
rect 11242 9072 11298 9081
rect 11152 9036 11204 9042
rect 11242 9007 11298 9016
rect 11152 8978 11204 8984
rect 11256 8906 11284 9007
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 10890 8732 11198 8741
rect 10890 8730 10896 8732
rect 10952 8730 10976 8732
rect 11032 8730 11056 8732
rect 11112 8730 11136 8732
rect 11192 8730 11198 8732
rect 10952 8678 10954 8730
rect 11134 8678 11136 8730
rect 10890 8676 10896 8678
rect 10952 8676 10976 8678
rect 11032 8676 11056 8678
rect 11112 8676 11136 8678
rect 11192 8676 11198 8678
rect 10890 8667 11198 8676
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 10890 7644 11198 7653
rect 10890 7642 10896 7644
rect 10952 7642 10976 7644
rect 11032 7642 11056 7644
rect 11112 7642 11136 7644
rect 11192 7642 11198 7644
rect 10952 7590 10954 7642
rect 11134 7590 11136 7642
rect 10890 7588 10896 7590
rect 10952 7588 10976 7590
rect 11032 7588 11056 7590
rect 11112 7588 11136 7590
rect 11192 7588 11198 7590
rect 10890 7579 11198 7588
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10704 3602 10732 4626
rect 10796 4010 10824 6870
rect 11256 6798 11284 7958
rect 11348 6866 11376 10134
rect 11440 10130 11468 11716
rect 11520 11698 11572 11704
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 8498 11468 9862
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 10890 6556 11198 6565
rect 10890 6554 10896 6556
rect 10952 6554 10976 6556
rect 11032 6554 11056 6556
rect 11112 6554 11136 6556
rect 11192 6554 11198 6556
rect 10952 6502 10954 6554
rect 11134 6502 11136 6554
rect 10890 6500 10896 6502
rect 10952 6500 10976 6502
rect 11032 6500 11056 6502
rect 11112 6500 11136 6502
rect 11192 6500 11198 6502
rect 10890 6491 11198 6500
rect 10890 5468 11198 5477
rect 10890 5466 10896 5468
rect 10952 5466 10976 5468
rect 11032 5466 11056 5468
rect 11112 5466 11136 5468
rect 11192 5466 11198 5468
rect 10952 5414 10954 5466
rect 11134 5414 11136 5466
rect 10890 5412 10896 5414
rect 10952 5412 10976 5414
rect 11032 5412 11056 5414
rect 11112 5412 11136 5414
rect 11192 5412 11198 5414
rect 10890 5403 11198 5412
rect 11256 5166 11284 6734
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 5914 11376 6598
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 10890 4380 11198 4389
rect 10890 4378 10896 4380
rect 10952 4378 10976 4380
rect 11032 4378 11056 4380
rect 11112 4378 11136 4380
rect 11192 4378 11198 4380
rect 10952 4326 10954 4378
rect 11134 4326 11136 4378
rect 10890 4324 10896 4326
rect 10952 4324 10976 4326
rect 11032 4324 11056 4326
rect 11112 4324 11136 4326
rect 11192 4324 11198 4326
rect 10890 4315 11198 4324
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 11072 3738 11100 4082
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11256 3602 11284 5102
rect 11348 4826 11376 5170
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 3738 11468 6054
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10890 3292 11198 3301
rect 10890 3290 10896 3292
rect 10952 3290 10976 3292
rect 11032 3290 11056 3292
rect 11112 3290 11136 3292
rect 11192 3290 11198 3292
rect 10952 3238 10954 3290
rect 11134 3238 11136 3290
rect 10890 3236 10896 3238
rect 10952 3236 10976 3238
rect 11032 3236 11056 3238
rect 11112 3236 11136 3238
rect 11192 3236 11198 3238
rect 10890 3227 11198 3236
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2650 10824 3130
rect 11256 3058 11284 3538
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11348 2854 11376 3334
rect 11532 2922 11560 11494
rect 11624 11218 11652 11562
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11624 10130 11652 10474
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9722 11744 9998
rect 11808 9908 11836 13942
rect 11886 12880 11942 12889
rect 11886 12815 11888 12824
rect 11940 12815 11942 12824
rect 11888 12786 11940 12792
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 12345 11928 12650
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11992 12209 12020 16050
rect 12084 13870 12112 16594
rect 12072 13864 12124 13870
rect 12070 13832 12072 13841
rect 12124 13832 12126 13841
rect 12268 13802 12296 17870
rect 12452 17338 12480 18294
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16590 12480 16934
rect 12440 16584 12492 16590
rect 12544 16561 12572 19858
rect 12728 19446 12756 20538
rect 12820 19786 12848 20538
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12624 19304 12676 19310
rect 12622 19272 12624 19281
rect 12676 19272 12678 19281
rect 12622 19207 12678 19216
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18426 12848 19178
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12440 16526 12492 16532
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 14074 12388 14214
rect 12544 14074 12572 16487
rect 12636 16454 12664 17138
rect 12820 16454 12848 17206
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12636 15706 12664 16118
rect 12820 16046 12848 16390
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12728 15706 12756 15982
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12070 13767 12126 13776
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12176 12730 12204 13670
rect 12360 13376 12388 13670
rect 12544 13530 12572 13874
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12268 13348 12388 13376
rect 12440 13388 12492 13394
rect 12268 13258 12296 13348
rect 12440 13330 12492 13336
rect 12452 13274 12480 13330
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12360 13246 12480 13274
rect 12360 12782 12388 13246
rect 12440 13184 12492 13190
rect 12728 13138 12756 13466
rect 12440 13126 12492 13132
rect 12452 13002 12480 13126
rect 12636 13110 12756 13138
rect 12636 13002 12664 13110
rect 12452 12974 12664 13002
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12348 12776 12400 12782
rect 12084 12434 12112 12718
rect 12176 12702 12296 12730
rect 12728 12753 12756 12786
rect 12714 12744 12770 12753
rect 12348 12718 12400 12724
rect 12164 12436 12216 12442
rect 12084 12406 12164 12434
rect 11978 12200 12034 12209
rect 11978 12135 12034 12144
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11900 11370 11928 11698
rect 11992 11540 12020 12135
rect 12084 11762 12112 12406
rect 12164 12378 12216 12384
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12176 11626 12204 12106
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 11992 11512 12112 11540
rect 11900 11342 12020 11370
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11900 10062 11928 10746
rect 11992 10606 12020 11342
rect 12084 10826 12112 11512
rect 12084 10798 12204 10826
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10198 12020 10542
rect 12084 10266 12112 10678
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11808 9880 11928 9908
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11610 9480 11666 9489
rect 11610 9415 11666 9424
rect 11624 7750 11652 9415
rect 11716 9110 11744 9658
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 6390 11652 7142
rect 11716 6848 11744 8298
rect 11808 7256 11836 9658
rect 11900 9518 11928 9880
rect 12176 9722 12204 10798
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9330 11928 9454
rect 12268 9330 12296 12702
rect 12636 12702 12714 12730
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12238 12480 12582
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12636 11286 12664 12702
rect 12714 12679 12770 12688
rect 12912 12434 12940 22170
rect 13004 20890 13032 25350
rect 13728 25298 13780 25304
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13188 24954 13216 25230
rect 13176 24948 13228 24954
rect 13176 24890 13228 24896
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13556 24410 13584 24686
rect 13740 24614 13768 25298
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13648 22438 13676 22510
rect 13636 22432 13688 22438
rect 13636 22374 13688 22380
rect 13648 22234 13676 22374
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13740 22030 13768 24550
rect 13832 23798 13860 25366
rect 14004 24880 14056 24886
rect 14004 24822 14056 24828
rect 14016 23866 14044 24822
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13820 23792 13872 23798
rect 14108 23746 14136 26250
rect 14844 26246 14872 28381
rect 15488 26382 15516 28381
rect 16417 26684 16725 26693
rect 16417 26682 16423 26684
rect 16479 26682 16503 26684
rect 16559 26682 16583 26684
rect 16639 26682 16663 26684
rect 16719 26682 16725 26684
rect 16479 26630 16481 26682
rect 16661 26630 16663 26682
rect 16417 26628 16423 26630
rect 16479 26628 16503 26630
rect 16559 26628 16583 26630
rect 16639 26628 16663 26630
rect 16719 26628 16725 26630
rect 16417 26619 16725 26628
rect 16776 26586 16804 28381
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 17420 26382 17448 28381
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14384 24954 14412 25162
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24206 14688 24550
rect 14648 24200 14700 24206
rect 14370 24168 14426 24177
rect 14648 24142 14700 24148
rect 14370 24103 14426 24112
rect 14384 24070 14412 24103
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 13820 23734 13872 23740
rect 14016 23718 14136 23746
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13096 21350 13124 21830
rect 13188 21690 13216 21830
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13648 21146 13676 21898
rect 13740 21622 13768 21966
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13740 21146 13768 21558
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20942 13860 21830
rect 13820 20936 13872 20942
rect 13004 20862 13124 20890
rect 13820 20878 13872 20884
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 20466 13032 20742
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12990 20088 13046 20097
rect 12990 20023 13046 20032
rect 13004 19378 13032 20023
rect 13096 19514 13124 20862
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13188 20602 13216 20810
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13096 19174 13124 19450
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13280 17882 13308 19450
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 15570 13216 16390
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13004 12850 13032 14010
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13280 12714 13308 12922
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 12820 12406 12940 12434
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 11900 9302 12020 9330
rect 11886 9208 11942 9217
rect 11886 9143 11942 9152
rect 11900 9042 11928 9143
rect 11992 9042 12020 9302
rect 12084 9302 12296 9330
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11900 8809 11928 8978
rect 11980 8832 12032 8838
rect 11886 8800 11942 8809
rect 11980 8774 12032 8780
rect 11886 8735 11942 8744
rect 11992 8498 12020 8774
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11900 7546 11928 7754
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12084 7342 12112 9302
rect 12360 9110 12388 9862
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12254 8800 12310 8809
rect 12254 8735 12310 8744
rect 12268 8566 12296 8735
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11888 7268 11940 7274
rect 11808 7228 11888 7256
rect 11888 7210 11940 7216
rect 11716 6820 11836 6848
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6458 11744 6666
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11808 3126 11836 6820
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6458 11928 6598
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 4622 12020 7278
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6186 12112 6802
rect 12176 6186 12204 8230
rect 12268 8022 12296 8366
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12452 7562 12480 10950
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12544 9897 12572 10474
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12544 9586 12572 9687
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12636 9489 12664 9930
rect 12728 9722 12756 9930
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12820 9568 12848 12406
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10305 12940 10406
rect 12898 10296 12954 10305
rect 12898 10231 12954 10240
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12912 9654 12940 9930
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12728 9540 12848 9568
rect 12622 9480 12678 9489
rect 12622 9415 12678 9424
rect 12636 8634 12664 9415
rect 12728 8922 12756 9540
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12728 8894 12848 8922
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8566 12756 8774
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12452 7546 12664 7562
rect 12452 7540 12676 7546
rect 12452 7534 12624 7540
rect 12624 7482 12676 7488
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12268 6866 12296 7278
rect 12452 7002 12480 7414
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4282 12020 4558
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12176 3194 12204 4694
rect 12268 4690 12296 6802
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 6458 12388 6666
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 5302 12480 5510
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12820 4842 12848 8894
rect 12912 8634 12940 8978
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12452 4814 12848 4842
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 12452 2514 12480 4814
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12728 4078 12756 4694
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12544 2650 12572 3402
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 10140 2440 10192 2446
rect 10416 2440 10468 2446
rect 10140 2382 10192 2388
rect 10336 2400 10416 2428
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 9048 800 9076 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10336 800 10364 2400
rect 11060 2440 11112 2446
rect 10416 2382 10468 2388
rect 10796 2400 11060 2428
rect 10796 1306 10824 2400
rect 11060 2382 11112 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 10890 2204 11198 2213
rect 10890 2202 10896 2204
rect 10952 2202 10976 2204
rect 11032 2202 11056 2204
rect 11112 2202 11136 2204
rect 11192 2202 11198 2204
rect 10952 2150 10954 2202
rect 11134 2150 11136 2202
rect 10890 2148 10896 2150
rect 10952 2148 10976 2150
rect 11032 2148 11056 2150
rect 11112 2148 11136 2150
rect 11192 2148 11198 2150
rect 10890 2139 11198 2148
rect 10796 1278 11008 1306
rect 10980 800 11008 1278
rect 12268 800 12296 2382
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12452 1698 12480 2246
rect 12636 1902 12664 3878
rect 12728 3398 12756 4014
rect 12912 4010 12940 4626
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 2038 12756 3334
rect 12806 2952 12862 2961
rect 12806 2887 12862 2896
rect 12820 2650 12848 2887
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 12624 1896 12676 1902
rect 12624 1838 12676 1844
rect 12440 1692 12492 1698
rect 12440 1634 12492 1640
rect 12912 800 12940 2246
rect 13004 1902 13032 12242
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13096 11286 13124 12106
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10130 13124 10406
rect 13280 10282 13308 12310
rect 13372 11218 13400 19654
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13924 18426 13952 18702
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13924 17882 13952 18362
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13464 15910 13492 16458
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12986 13492 13262
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13556 10674 13584 14826
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 13394 13676 14282
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12986 13676 13330
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13648 12442 13676 12786
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13740 12238 13768 17478
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16697 13860 17070
rect 13818 16688 13874 16697
rect 13818 16623 13874 16632
rect 14016 14385 14044 23718
rect 14476 23322 14504 24006
rect 14554 23760 14610 23769
rect 14660 23746 14688 24142
rect 14610 23718 14780 23746
rect 14554 23695 14610 23704
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22234 14136 22918
rect 14292 22778 14320 23054
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14200 22506 14228 22714
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14476 21978 14504 23258
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14568 22574 14596 23054
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14384 21950 14504 21978
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 20942 14228 21422
rect 14384 20942 14412 21950
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14476 20942 14504 21830
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14200 19378 14228 19994
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 18970 14228 19314
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 15910 14228 16390
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 14408 14148 14414
rect 14002 14376 14058 14385
rect 14096 14350 14148 14356
rect 14002 14311 14058 14320
rect 14108 13326 14136 14350
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 14200 11354 14228 15846
rect 14292 14618 14320 20742
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18290 14412 19246
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14476 17610 14504 18906
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14568 16726 14596 22510
rect 14752 20942 14780 23718
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14660 20058 14688 20878
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14646 19000 14702 19009
rect 14752 18970 14780 19178
rect 14646 18935 14702 18944
rect 14740 18964 14792 18970
rect 14660 18766 14688 18935
rect 14740 18906 14792 18912
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14738 18728 14794 18737
rect 14738 18663 14740 18672
rect 14792 18663 14794 18672
rect 14740 18634 14792 18640
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14568 15570 14596 16662
rect 14660 16590 14688 18294
rect 14844 17746 14872 19382
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14936 18698 14964 19110
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14752 17338 14780 17682
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 15028 17218 15056 26250
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15120 24682 15148 25094
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15212 21593 15240 26250
rect 16212 26036 16264 26042
rect 16212 25978 16264 25984
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15842 25800 15898 25809
rect 15842 25735 15898 25744
rect 15856 25498 15884 25735
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15304 24206 15332 24890
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15488 24070 15516 24754
rect 15580 24410 15608 24754
rect 15856 24698 15884 25434
rect 15764 24670 15884 24698
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15672 23866 15700 24142
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15672 23322 15700 23666
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15672 22166 15700 22646
rect 15764 22574 15792 24670
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 24410 15884 24550
rect 15948 24410 15976 25842
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15948 23866 15976 24346
rect 16132 24206 16160 25774
rect 16224 24750 16252 25978
rect 16417 25596 16725 25605
rect 16417 25594 16423 25596
rect 16479 25594 16503 25596
rect 16559 25594 16583 25596
rect 16639 25594 16663 25596
rect 16719 25594 16725 25596
rect 16479 25542 16481 25594
rect 16661 25542 16663 25594
rect 16417 25540 16423 25542
rect 16479 25540 16503 25542
rect 16559 25540 16583 25542
rect 16639 25540 16663 25542
rect 16719 25540 16725 25542
rect 16417 25531 16725 25540
rect 16868 25498 16896 26250
rect 17077 26140 17385 26149
rect 17077 26138 17083 26140
rect 17139 26138 17163 26140
rect 17219 26138 17243 26140
rect 17299 26138 17323 26140
rect 17379 26138 17385 26140
rect 17139 26086 17141 26138
rect 17321 26086 17323 26138
rect 17077 26084 17083 26086
rect 17139 26084 17163 26086
rect 17219 26084 17243 26086
rect 17299 26084 17323 26086
rect 17379 26084 17385 26086
rect 17077 26075 17385 26084
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 16672 25288 16724 25294
rect 16868 25242 16896 25434
rect 16724 25236 16896 25242
rect 16672 25230 16896 25236
rect 16684 25214 16896 25230
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24954 16620 25094
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16684 24682 16712 25214
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16868 24886 16896 25094
rect 16856 24880 16908 24886
rect 16856 24822 16908 24828
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16672 24676 16724 24682
rect 16672 24618 16724 24624
rect 16417 24508 16725 24517
rect 16417 24506 16423 24508
rect 16479 24506 16503 24508
rect 16559 24506 16583 24508
rect 16639 24506 16663 24508
rect 16719 24506 16725 24508
rect 16479 24454 16481 24506
rect 16661 24454 16663 24506
rect 16417 24452 16423 24454
rect 16479 24452 16503 24454
rect 16559 24452 16583 24454
rect 16639 24452 16663 24454
rect 16719 24452 16725 24454
rect 16417 24443 16725 24452
rect 16394 24304 16450 24313
rect 16394 24239 16450 24248
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16028 23724 16080 23730
rect 15948 23684 16028 23712
rect 15948 23322 15976 23684
rect 16028 23666 16080 23672
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15948 22234 15976 22578
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15198 21584 15254 21593
rect 15198 21519 15254 21528
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 20058 15424 20266
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15106 19952 15162 19961
rect 15106 19887 15108 19896
rect 15160 19887 15162 19896
rect 15108 19858 15160 19864
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15396 19718 15424 19790
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15384 19372 15436 19378
rect 15304 19320 15384 19334
rect 15304 19314 15436 19320
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15304 19306 15424 19314
rect 15120 18766 15148 19246
rect 15212 18850 15240 19246
rect 15304 18970 15332 19306
rect 15488 19292 15516 21354
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15580 19446 15608 19790
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15672 19310 15700 22102
rect 15936 20460 15988 20466
rect 16040 20448 16068 23530
rect 16224 23254 16252 24006
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 20534 16160 23054
rect 16224 22574 16252 23190
rect 16316 23118 16344 23802
rect 16408 23594 16436 24239
rect 16776 23798 16804 24754
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16764 23792 16816 23798
rect 16764 23734 16816 23740
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16417 23420 16725 23429
rect 16417 23418 16423 23420
rect 16479 23418 16503 23420
rect 16559 23418 16583 23420
rect 16639 23418 16663 23420
rect 16719 23418 16725 23420
rect 16479 23366 16481 23418
rect 16661 23366 16663 23418
rect 16417 23364 16423 23366
rect 16479 23364 16503 23366
rect 16559 23364 16583 23366
rect 16639 23364 16663 23366
rect 16719 23364 16725 23366
rect 16417 23355 16725 23364
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 22030 16252 22374
rect 16316 22234 16344 22918
rect 16417 22332 16725 22341
rect 16417 22330 16423 22332
rect 16479 22330 16503 22332
rect 16559 22330 16583 22332
rect 16639 22330 16663 22332
rect 16719 22330 16725 22332
rect 16479 22278 16481 22330
rect 16661 22278 16663 22330
rect 16417 22276 16423 22278
rect 16479 22276 16503 22278
rect 16559 22276 16583 22278
rect 16639 22276 16663 22278
rect 16719 22276 16725 22278
rect 16417 22267 16725 22276
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16776 22094 16804 23054
rect 16868 22760 16896 24346
rect 16960 24274 16988 25094
rect 17077 25052 17385 25061
rect 17077 25050 17083 25052
rect 17139 25050 17163 25052
rect 17219 25050 17243 25052
rect 17299 25050 17323 25052
rect 17379 25050 17385 25052
rect 17139 24998 17141 25050
rect 17321 24998 17323 25050
rect 17077 24996 17083 24998
rect 17139 24996 17163 24998
rect 17219 24996 17243 24998
rect 17299 24996 17323 24998
rect 17379 24996 17385 24998
rect 17077 24987 17385 24996
rect 17420 24954 17448 25434
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 24426 17356 24686
rect 17052 24398 17356 24426
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17052 24154 17080 24398
rect 17132 24336 17184 24342
rect 17420 24290 17448 24890
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 17184 24284 17448 24290
rect 17132 24278 17448 24284
rect 17144 24262 17448 24278
rect 17604 24290 17632 24822
rect 17696 24426 17724 26522
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17788 25498 17816 25842
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17880 25362 17908 25774
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17788 24886 17816 25094
rect 17776 24880 17828 24886
rect 17776 24822 17828 24828
rect 17696 24398 17908 24426
rect 17604 24262 17724 24290
rect 17420 24206 17448 24262
rect 17132 24200 17184 24206
rect 17052 24148 17132 24154
rect 17052 24142 17184 24148
rect 17408 24200 17460 24206
rect 17500 24200 17552 24206
rect 17408 24142 17460 24148
rect 17498 24168 17500 24177
rect 17552 24168 17554 24177
rect 17052 24126 17172 24142
rect 17498 24103 17554 24112
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23526 16988 24006
rect 17077 23964 17385 23973
rect 17077 23962 17083 23964
rect 17139 23962 17163 23964
rect 17219 23962 17243 23964
rect 17299 23962 17323 23964
rect 17379 23962 17385 23964
rect 17139 23910 17141 23962
rect 17321 23910 17323 23962
rect 17077 23908 17083 23910
rect 17139 23908 17163 23910
rect 17219 23908 17243 23910
rect 17299 23908 17323 23910
rect 17379 23908 17385 23910
rect 17077 23899 17385 23908
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16960 23322 16988 23462
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17077 22876 17385 22885
rect 17077 22874 17083 22876
rect 17139 22874 17163 22876
rect 17219 22874 17243 22876
rect 17299 22874 17323 22876
rect 17379 22874 17385 22876
rect 17139 22822 17141 22874
rect 17321 22822 17323 22874
rect 17077 22820 17083 22822
rect 17139 22820 17163 22822
rect 17219 22820 17243 22822
rect 17299 22820 17323 22822
rect 17379 22820 17385 22822
rect 17077 22811 17385 22820
rect 17420 22778 17448 23054
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17316 22772 17368 22778
rect 16868 22732 17080 22760
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16684 22066 16804 22094
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16224 21690 16252 21966
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16684 21622 16712 22066
rect 16960 22030 16988 22374
rect 17052 22098 17080 22732
rect 17316 22714 17368 22720
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17328 22574 17356 22714
rect 17512 22710 17540 22918
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17604 22574 17632 23666
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17328 22234 17356 22510
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17420 22030 17448 22442
rect 17696 22386 17724 24262
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17604 22358 17724 22386
rect 17604 22137 17632 22358
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17590 22128 17646 22137
rect 17590 22063 17646 22072
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 16776 21690 16804 21966
rect 16856 21888 16908 21894
rect 17144 21876 17172 21966
rect 16856 21830 16908 21836
rect 16960 21848 17172 21876
rect 17500 21888 17552 21894
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16417 21244 16725 21253
rect 16417 21242 16423 21244
rect 16479 21242 16503 21244
rect 16559 21242 16583 21244
rect 16639 21242 16663 21244
rect 16719 21242 16725 21244
rect 16479 21190 16481 21242
rect 16661 21190 16663 21242
rect 16417 21188 16423 21190
rect 16479 21188 16503 21190
rect 16559 21188 16583 21190
rect 16639 21188 16663 21190
rect 16719 21188 16725 21190
rect 16417 21179 16725 21188
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 15988 20420 16068 20448
rect 15936 20402 15988 20408
rect 15948 20330 15976 20402
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 16132 19990 16160 20470
rect 16120 19984 16172 19990
rect 16120 19926 16172 19932
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15660 19304 15712 19310
rect 15488 19264 15608 19292
rect 15488 19174 15516 19264
rect 15476 19168 15528 19174
rect 15580 19156 15608 19264
rect 15660 19246 15712 19252
rect 15764 19224 15792 19790
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15844 19236 15896 19242
rect 15764 19196 15844 19224
rect 15844 19178 15896 19184
rect 15580 19128 15700 19156
rect 15476 19110 15528 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15476 18896 15528 18902
rect 15212 18822 15332 18850
rect 15476 18838 15528 18844
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15120 18630 15148 18702
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 15106 18320 15162 18329
rect 15212 18290 15240 18702
rect 15106 18255 15108 18264
rect 15160 18255 15162 18264
rect 15200 18284 15252 18290
rect 15108 18226 15160 18232
rect 15200 18226 15252 18232
rect 15028 17190 15148 17218
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14936 16658 14964 16934
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 13258 14320 13670
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 12238 14504 12718
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 13740 10674 13768 11290
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13924 11121 13952 11222
rect 14568 11150 14596 15506
rect 15028 15094 15056 16390
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 13938 14780 14894
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 12918 14872 13806
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14936 12714 14964 13738
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 15120 12434 15148 17190
rect 15304 17134 15332 18822
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15396 18358 15424 18634
rect 15488 18358 15516 18838
rect 15568 18760 15620 18766
rect 15672 18737 15700 19128
rect 15842 19000 15898 19009
rect 15948 18970 15976 19246
rect 15842 18935 15844 18944
rect 15896 18935 15898 18944
rect 15936 18964 15988 18970
rect 15844 18906 15896 18912
rect 16040 18952 16068 19654
rect 16132 19378 16160 19790
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16040 18924 16160 18952
rect 15936 18906 15988 18912
rect 15844 18828 15896 18834
rect 16132 18816 16160 18924
rect 15844 18770 15896 18776
rect 16040 18788 16160 18816
rect 15752 18760 15804 18766
rect 15568 18702 15620 18708
rect 15658 18728 15714 18737
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15580 18290 15608 18702
rect 15752 18702 15804 18708
rect 15658 18663 15714 18672
rect 15672 18306 15700 18663
rect 15764 18426 15792 18702
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15856 18358 15884 18770
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18352 15896 18358
rect 15568 18284 15620 18290
rect 15672 18278 15792 18306
rect 15844 18294 15896 18300
rect 15568 18226 15620 18232
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 17610 15424 18022
rect 15580 17882 15608 18226
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 17202 15424 17546
rect 15488 17202 15516 17682
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16046 15332 17070
rect 15396 16522 15424 17138
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15488 16182 15516 17138
rect 15580 16998 15608 17206
rect 15672 16998 15700 17274
rect 15764 17202 15792 18278
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15856 17270 15884 18090
rect 15948 17882 15976 18362
rect 16040 18290 16068 18788
rect 16224 18340 16252 20878
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 20058 16344 20402
rect 16417 20156 16725 20165
rect 16417 20154 16423 20156
rect 16479 20154 16503 20156
rect 16559 20154 16583 20156
rect 16639 20154 16663 20156
rect 16719 20154 16725 20156
rect 16479 20102 16481 20154
rect 16661 20102 16663 20154
rect 16417 20100 16423 20102
rect 16479 20100 16503 20102
rect 16559 20100 16583 20102
rect 16639 20100 16663 20102
rect 16719 20100 16725 20102
rect 16417 20091 16725 20100
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16316 19922 16344 19994
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16592 19446 16620 19722
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16316 18970 16344 19314
rect 16684 19174 16712 19314
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16417 19068 16725 19077
rect 16417 19066 16423 19068
rect 16479 19066 16503 19068
rect 16559 19066 16583 19068
rect 16639 19066 16663 19068
rect 16719 19066 16725 19068
rect 16479 19014 16481 19066
rect 16661 19014 16663 19066
rect 16417 19012 16423 19014
rect 16479 19012 16503 19014
rect 16559 19012 16583 19014
rect 16639 19012 16663 19014
rect 16719 19012 16725 19014
rect 16417 19003 16725 19012
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16776 18766 16804 19110
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16500 18426 16528 18702
rect 16684 18426 16712 18702
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16396 18352 16448 18358
rect 16224 18312 16396 18340
rect 16684 18329 16712 18362
rect 16396 18294 16448 18300
rect 16670 18320 16726 18329
rect 16028 18284 16080 18290
rect 16670 18255 16726 18264
rect 16028 18226 16080 18232
rect 16684 18068 16712 18255
rect 16776 18222 16804 18702
rect 16868 18698 16896 21830
rect 16960 21554 16988 21848
rect 17500 21830 17552 21836
rect 17077 21788 17385 21797
rect 17077 21786 17083 21788
rect 17139 21786 17163 21788
rect 17219 21786 17243 21788
rect 17299 21786 17323 21788
rect 17379 21786 17385 21788
rect 17139 21734 17141 21786
rect 17321 21734 17323 21786
rect 17077 21732 17083 21734
rect 17139 21732 17163 21734
rect 17219 21732 17243 21734
rect 17299 21732 17323 21734
rect 17379 21732 17385 21734
rect 17077 21723 17385 21732
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 16948 21412 17000 21418
rect 17236 21400 17264 21490
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17000 21372 17264 21400
rect 16948 21354 17000 21360
rect 17420 20806 17448 21422
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17077 20700 17385 20709
rect 17077 20698 17083 20700
rect 17139 20698 17163 20700
rect 17219 20698 17243 20700
rect 17299 20698 17323 20700
rect 17379 20698 17385 20700
rect 17139 20646 17141 20698
rect 17321 20646 17323 20698
rect 17077 20644 17083 20646
rect 17139 20644 17163 20646
rect 17219 20644 17243 20646
rect 17299 20644 17323 20646
rect 17379 20644 17385 20646
rect 17077 20635 17385 20644
rect 17512 20058 17540 21830
rect 17604 21418 17632 21966
rect 17696 21418 17724 22170
rect 17788 22030 17816 22578
rect 17880 22234 17908 24398
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17866 21992 17922 22001
rect 17866 21927 17922 21936
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17684 21412 17736 21418
rect 17684 21354 17736 21360
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17077 19612 17385 19621
rect 17077 19610 17083 19612
rect 17139 19610 17163 19612
rect 17219 19610 17243 19612
rect 17299 19610 17323 19612
rect 17379 19610 17385 19612
rect 17139 19558 17141 19610
rect 17321 19558 17323 19610
rect 17077 19556 17083 19558
rect 17139 19556 17163 19558
rect 17219 19556 17243 19558
rect 17299 19556 17323 19558
rect 17379 19556 17385 19558
rect 17077 19547 17385 19556
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 17052 18630 17080 19382
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17077 18524 17385 18533
rect 17077 18522 17083 18524
rect 17139 18522 17163 18524
rect 17219 18522 17243 18524
rect 17299 18522 17323 18524
rect 17379 18522 17385 18524
rect 17139 18470 17141 18522
rect 17321 18470 17323 18522
rect 17077 18468 17083 18470
rect 17139 18468 17163 18470
rect 17219 18468 17243 18470
rect 17299 18468 17323 18470
rect 17379 18468 17385 18470
rect 17077 18459 17385 18468
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 17052 18170 17080 18226
rect 17052 18142 17172 18170
rect 17144 18086 17172 18142
rect 17040 18080 17092 18086
rect 16684 18040 16804 18068
rect 16417 17980 16725 17989
rect 16417 17978 16423 17980
rect 16479 17978 16503 17980
rect 16559 17978 16583 17980
rect 16639 17978 16663 17980
rect 16719 17978 16725 17980
rect 16479 17926 16481 17978
rect 16661 17926 16663 17978
rect 16417 17924 16423 17926
rect 16479 17924 16503 17926
rect 16559 17924 16583 17926
rect 16639 17924 16663 17926
rect 16719 17924 16725 17926
rect 16417 17915 16725 17924
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16040 17270 16068 17478
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15580 16658 15608 16934
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15764 16250 15792 16594
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 15570 15332 15846
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15200 15088 15252 15094
rect 15198 15056 15200 15065
rect 15252 15056 15254 15065
rect 15396 15026 15424 15302
rect 15198 14991 15254 15000
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14482 15516 14894
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 12918 15240 14214
rect 15580 14074 15608 14282
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 12918 15332 13874
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15028 12406 15148 12434
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14556 11144 14608 11150
rect 13910 11112 13966 11121
rect 14556 11086 14608 11092
rect 13910 11047 13966 11056
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10470 13768 10610
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13176 10260 13228 10266
rect 13280 10254 13400 10282
rect 13176 10202 13228 10208
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9382 13124 10066
rect 13188 10062 13216 10202
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13188 9722 13216 9998
rect 13280 9761 13308 10134
rect 13266 9752 13322 9761
rect 13176 9716 13228 9722
rect 13266 9687 13322 9696
rect 13176 9658 13228 9664
rect 13280 9654 13308 9687
rect 13268 9648 13320 9654
rect 13174 9616 13230 9625
rect 13268 9590 13320 9596
rect 13174 9551 13230 9560
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13188 9178 13216 9551
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13372 8022 13400 10254
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9489 13492 9998
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13648 9586 13676 9930
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13450 9480 13506 9489
rect 13450 9415 13506 9424
rect 13556 9217 13584 9522
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13542 9072 13598 9081
rect 13542 9007 13598 9016
rect 13556 8974 13584 9007
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13832 8090 13860 8434
rect 13924 8090 13952 11047
rect 14752 11014 14780 11290
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14016 9110 14044 10678
rect 14292 10062 14320 10950
rect 14556 10464 14608 10470
rect 14608 10424 14688 10452
rect 14556 10406 14608 10412
rect 14660 10062 14688 10424
rect 14752 10130 14780 10950
rect 14830 10296 14886 10305
rect 14830 10231 14886 10240
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14844 9926 14872 10231
rect 14936 10198 14964 10950
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14108 9586 14136 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14188 9376 14240 9382
rect 14292 9353 14320 9454
rect 14188 9318 14240 9324
rect 14278 9344 14334 9353
rect 14200 9178 14228 9318
rect 14278 9279 14334 9288
rect 14844 9178 14872 9454
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4690 13308 4966
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13372 3670 13400 7958
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 3194 13308 3334
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 13280 1562 13308 2790
rect 13464 1834 13492 7210
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5642 13676 6054
rect 13924 5914 13952 6122
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13740 4010 13768 5646
rect 14016 5370 14044 9046
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8634 14228 8774
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14108 6390 14136 7414
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13832 4826 13860 5170
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 4146 13952 4422
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13648 2774 13676 3606
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13648 2746 13768 2774
rect 13740 2530 13768 2746
rect 13832 2650 13860 3334
rect 13924 3058 13952 3334
rect 14108 3126 14136 4966
rect 14200 3670 14228 7686
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14292 5642 14320 6938
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14384 5710 14412 6122
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14292 4758 14320 5578
rect 14476 5273 14504 8910
rect 14844 6458 14872 9114
rect 15028 8378 15056 12406
rect 15212 9994 15240 12718
rect 15396 12442 15424 13194
rect 15764 12782 15792 15982
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 15570 15976 15846
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16132 15434 16160 17478
rect 16224 17338 16252 17614
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 16182 16252 16526
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16224 15910 16252 16118
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16316 15722 16344 17614
rect 16417 16892 16725 16901
rect 16417 16890 16423 16892
rect 16479 16890 16503 16892
rect 16559 16890 16583 16892
rect 16639 16890 16663 16892
rect 16719 16890 16725 16892
rect 16479 16838 16481 16890
rect 16661 16838 16663 16890
rect 16417 16836 16423 16838
rect 16479 16836 16503 16838
rect 16559 16836 16583 16838
rect 16639 16836 16663 16838
rect 16719 16836 16725 16838
rect 16417 16827 16725 16836
rect 16417 15804 16725 15813
rect 16417 15802 16423 15804
rect 16479 15802 16503 15804
rect 16559 15802 16583 15804
rect 16639 15802 16663 15804
rect 16719 15802 16725 15804
rect 16479 15750 16481 15802
rect 16661 15750 16663 15802
rect 16417 15748 16423 15750
rect 16479 15748 16503 15750
rect 16559 15748 16583 15750
rect 16639 15748 16663 15750
rect 16719 15748 16725 15750
rect 16417 15739 16725 15748
rect 16224 15694 16344 15722
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 16224 15094 16252 15694
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15752 12776 15804 12782
rect 15856 12753 15884 13126
rect 16132 12986 16160 13874
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15752 12718 15804 12724
rect 15842 12744 15898 12753
rect 15842 12679 15898 12688
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10062 15332 10542
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 8906 15148 9318
rect 15212 9110 15240 9930
rect 15304 9518 15332 9998
rect 15396 9654 15424 11698
rect 15580 10418 15608 11698
rect 15856 11665 15884 12679
rect 16040 12434 16068 12854
rect 16040 12406 16160 12434
rect 15842 11656 15898 11665
rect 15842 11591 15898 11600
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11218 15884 11494
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15488 10390 15608 10418
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15488 9450 15516 10390
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15580 9602 15608 10134
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15672 9926 15700 9998
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15580 9586 15700 9602
rect 15580 9580 15712 9586
rect 15580 9574 15660 9580
rect 15660 9522 15712 9528
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15028 8350 15148 8378
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 7818 15056 8230
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15120 7274 15148 8350
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 7002 15056 7142
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15396 6934 15424 7210
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15016 6180 15068 6186
rect 14936 6140 15016 6168
rect 14832 6112 14884 6118
rect 14936 6100 14964 6140
rect 15016 6122 15068 6128
rect 14884 6072 14964 6100
rect 14832 6054 14884 6060
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14462 5264 14518 5273
rect 14462 5199 14464 5208
rect 14516 5199 14518 5208
rect 14464 5170 14516 5176
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14292 4282 14320 4694
rect 14660 4690 14688 5714
rect 14844 5234 14872 6054
rect 15304 5914 15332 6258
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15212 5794 15240 5850
rect 15212 5766 15424 5794
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5234 15332 5578
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14752 4282 14780 5102
rect 14844 4282 14872 5170
rect 15396 5148 15424 5766
rect 15488 5352 15516 9386
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15672 8634 15700 8842
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7546 15608 7754
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15672 7410 15700 8570
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15672 6458 15700 6666
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6361 15792 11086
rect 16132 10674 16160 12406
rect 16224 11218 16252 15030
rect 16316 14074 16344 15370
rect 16417 14716 16725 14725
rect 16417 14714 16423 14716
rect 16479 14714 16503 14716
rect 16559 14714 16583 14716
rect 16639 14714 16663 14716
rect 16719 14714 16725 14716
rect 16479 14662 16481 14714
rect 16661 14662 16663 14714
rect 16417 14660 16423 14662
rect 16479 14660 16503 14662
rect 16559 14660 16583 14662
rect 16639 14660 16663 14662
rect 16719 14660 16725 14662
rect 16417 14651 16725 14660
rect 16672 14476 16724 14482
rect 16776 14464 16804 18040
rect 17040 18022 17092 18028
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17052 17678 17080 18022
rect 17328 17814 17356 18022
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17077 17436 17385 17445
rect 17077 17434 17083 17436
rect 17139 17434 17163 17436
rect 17219 17434 17243 17436
rect 17299 17434 17323 17436
rect 17379 17434 17385 17436
rect 17139 17382 17141 17434
rect 17321 17382 17323 17434
rect 17077 17380 17083 17382
rect 17139 17380 17163 17382
rect 17219 17380 17243 17382
rect 17299 17380 17323 17382
rect 17379 17380 17385 17382
rect 17077 17371 17385 17380
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16868 16726 16896 17070
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16960 15366 16988 16730
rect 17077 16348 17385 16357
rect 17077 16346 17083 16348
rect 17139 16346 17163 16348
rect 17219 16346 17243 16348
rect 17299 16346 17323 16348
rect 17379 16346 17385 16348
rect 17139 16294 17141 16346
rect 17321 16294 17323 16346
rect 17077 16292 17083 16294
rect 17139 16292 17163 16294
rect 17219 16292 17243 16294
rect 17299 16292 17323 16294
rect 17379 16292 17385 16294
rect 17077 16283 17385 16292
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17077 15260 17385 15269
rect 17077 15258 17083 15260
rect 17139 15258 17163 15260
rect 17219 15258 17243 15260
rect 17299 15258 17323 15260
rect 17379 15258 17385 15260
rect 17139 15206 17141 15258
rect 17321 15206 17323 15258
rect 17077 15204 17083 15206
rect 17139 15204 17163 15206
rect 17219 15204 17243 15206
rect 17299 15204 17323 15206
rect 17379 15204 17385 15206
rect 17077 15195 17385 15204
rect 17420 15162 17448 18294
rect 17512 18290 17540 18702
rect 17604 18630 17632 21354
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17788 18290 17816 18634
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17788 18154 17816 18226
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 16250 17816 16390
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17512 15892 17540 16186
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17604 16046 17632 16118
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17512 15864 17632 15892
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 16724 14436 16804 14464
rect 16672 14418 16724 14424
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16684 13938 16712 14418
rect 17077 14172 17385 14181
rect 17077 14170 17083 14172
rect 17139 14170 17163 14172
rect 17219 14170 17243 14172
rect 17299 14170 17323 14172
rect 17379 14170 17385 14172
rect 17139 14118 17141 14170
rect 17321 14118 17323 14170
rect 17077 14116 17083 14118
rect 17139 14116 17163 14118
rect 17219 14116 17243 14118
rect 17299 14116 17323 14118
rect 17379 14116 17385 14118
rect 17077 14107 17385 14116
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16417 13628 16725 13637
rect 16417 13626 16423 13628
rect 16479 13626 16503 13628
rect 16559 13626 16583 13628
rect 16639 13626 16663 13628
rect 16719 13626 16725 13628
rect 16479 13574 16481 13626
rect 16661 13574 16663 13626
rect 16417 13572 16423 13574
rect 16479 13572 16503 13574
rect 16559 13572 16583 13574
rect 16639 13572 16663 13574
rect 16719 13572 16725 13574
rect 16417 13563 16725 13572
rect 16776 13530 16804 13670
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16578 13424 16634 13433
rect 16684 13410 16712 13466
rect 16868 13410 16896 13738
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16684 13382 16896 13410
rect 16578 13359 16634 13368
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12986 16344 13262
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16592 12918 16620 13359
rect 17420 13258 17448 13670
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17077 13084 17385 13093
rect 17077 13082 17083 13084
rect 17139 13082 17163 13084
rect 17219 13082 17243 13084
rect 17299 13082 17323 13084
rect 17379 13082 17385 13084
rect 17139 13030 17141 13082
rect 17321 13030 17323 13082
rect 17077 13028 17083 13030
rect 17139 13028 17163 13030
rect 17219 13028 17243 13030
rect 17299 13028 17323 13030
rect 17379 13028 17385 13030
rect 17077 13019 17385 13028
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 17408 12844 17460 12850
rect 17512 12832 17540 15574
rect 17604 15434 17632 15864
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17460 12804 17540 12832
rect 17408 12786 17460 12792
rect 17132 12776 17184 12782
rect 16960 12736 17132 12764
rect 16417 12540 16725 12549
rect 16417 12538 16423 12540
rect 16479 12538 16503 12540
rect 16559 12538 16583 12540
rect 16639 12538 16663 12540
rect 16719 12538 16725 12540
rect 16479 12486 16481 12538
rect 16661 12486 16663 12538
rect 16417 12484 16423 12486
rect 16479 12484 16503 12486
rect 16559 12484 16583 12486
rect 16639 12484 16663 12486
rect 16719 12484 16725 12486
rect 16417 12475 16725 12484
rect 16417 11452 16725 11461
rect 16417 11450 16423 11452
rect 16479 11450 16503 11452
rect 16559 11450 16583 11452
rect 16639 11450 16663 11452
rect 16719 11450 16725 11452
rect 16479 11398 16481 11450
rect 16661 11398 16663 11450
rect 16417 11396 16423 11398
rect 16479 11396 16503 11398
rect 16559 11396 16583 11398
rect 16639 11396 16663 11398
rect 16719 11396 16725 11398
rect 16417 11387 16725 11396
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15856 10538 15884 10610
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 16040 10266 16068 10610
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16132 10010 16160 10610
rect 16500 10538 16528 10950
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10146 16252 10406
rect 16316 10248 16344 10474
rect 16417 10364 16725 10373
rect 16417 10362 16423 10364
rect 16479 10362 16503 10364
rect 16559 10362 16583 10364
rect 16639 10362 16663 10364
rect 16719 10362 16725 10364
rect 16479 10310 16481 10362
rect 16661 10310 16663 10362
rect 16417 10308 16423 10310
rect 16479 10308 16503 10310
rect 16559 10308 16583 10310
rect 16639 10308 16663 10310
rect 16719 10308 16725 10310
rect 16417 10299 16725 10308
rect 16316 10220 16620 10248
rect 16224 10118 16344 10146
rect 16132 9982 16252 10010
rect 15844 9920 15896 9926
rect 16120 9920 16172 9926
rect 15844 9862 15896 9868
rect 16040 9880 16120 9908
rect 15856 9586 15884 9862
rect 16040 9586 16068 9880
rect 16120 9862 16172 9868
rect 16224 9674 16252 9982
rect 16132 9646 16252 9674
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15856 9450 15884 9522
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 16040 9178 16068 9522
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16028 8968 16080 8974
rect 16132 8956 16160 9646
rect 16080 8928 16160 8956
rect 16212 8968 16264 8974
rect 16028 8910 16080 8916
rect 16212 8910 16264 8916
rect 16224 8090 16252 8910
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16224 7478 16252 8026
rect 16212 7472 16264 7478
rect 16212 7414 16264 7420
rect 16316 7342 16344 10118
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9994 16528 10066
rect 16488 9988 16540 9994
rect 16592 9976 16620 10220
rect 16776 10044 16804 11018
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16868 10266 16896 10474
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16856 10056 16908 10062
rect 16776 10016 16856 10044
rect 16856 9998 16908 10004
rect 16592 9948 16804 9976
rect 16488 9930 16540 9936
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9761 16436 9862
rect 16394 9752 16450 9761
rect 16394 9687 16450 9696
rect 16500 9586 16528 9930
rect 16578 9888 16634 9897
rect 16578 9823 16634 9832
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16592 9518 16620 9823
rect 16670 9752 16726 9761
rect 16670 9687 16726 9696
rect 16776 9704 16804 9948
rect 16960 9897 16988 12736
rect 17132 12718 17184 12724
rect 17420 12306 17448 12786
rect 17604 12764 17632 15370
rect 17880 15178 17908 21927
rect 17788 15150 17908 15178
rect 17788 13802 17816 15150
rect 17972 15026 18000 26386
rect 18064 26382 18092 28381
rect 19076 26586 19104 28478
rect 19982 28381 20038 29181
rect 20626 28381 20682 29181
rect 21270 28381 21326 29181
rect 21914 28506 21970 29181
rect 22926 28656 22982 28665
rect 22926 28591 22982 28600
rect 21914 28478 22048 28506
rect 21914 28381 21970 28478
rect 19996 26586 20024 28381
rect 20640 26602 20668 28381
rect 20640 26586 20760 26602
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 19984 26580 20036 26586
rect 20640 26580 20772 26586
rect 20640 26574 20720 26580
rect 19984 26522 20036 26528
rect 20720 26522 20772 26528
rect 18236 26512 18288 26518
rect 18236 26454 18288 26460
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18248 25294 18276 26454
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18524 25401 18552 25638
rect 18800 25498 18828 25910
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 18510 25392 18566 25401
rect 18510 25327 18512 25336
rect 18564 25327 18566 25336
rect 18512 25298 18564 25304
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18156 24682 18184 24754
rect 19352 24750 19380 25230
rect 19444 24954 19472 26250
rect 21284 26246 21312 28381
rect 22020 26466 22048 28478
rect 22604 26684 22912 26693
rect 22604 26682 22610 26684
rect 22666 26682 22690 26684
rect 22746 26682 22770 26684
rect 22826 26682 22850 26684
rect 22906 26682 22912 26684
rect 22666 26630 22668 26682
rect 22848 26630 22850 26682
rect 22604 26628 22610 26630
rect 22666 26628 22690 26630
rect 22746 26628 22770 26630
rect 22826 26628 22850 26630
rect 22906 26628 22912 26630
rect 22604 26619 22912 26628
rect 22836 26512 22888 26518
rect 22020 26438 22140 26466
rect 22836 26454 22888 26460
rect 22112 26382 22140 26438
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 21732 26308 21784 26314
rect 21732 26250 21784 26256
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 19708 25832 19760 25838
rect 19708 25774 19760 25780
rect 19720 25498 19748 25774
rect 20364 25498 20392 25842
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 20352 25492 20404 25498
rect 20352 25434 20404 25440
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18248 24138 18276 24550
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 19352 23798 19380 24686
rect 19536 24206 19564 25162
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19628 23866 19656 24686
rect 19800 24608 19852 24614
rect 19852 24568 19932 24596
rect 19800 24550 19852 24556
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19352 22642 19380 23734
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19536 23254 19564 23530
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19720 22778 19748 22918
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 21486 18092 22374
rect 19248 22094 19300 22098
rect 19352 22094 19380 22578
rect 19248 22092 19380 22094
rect 19300 22066 19380 22092
rect 19248 22034 19300 22040
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18340 21554 18368 21830
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18878 20360 18934 20369
rect 18340 20058 18368 20334
rect 18878 20295 18934 20304
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19446 18092 19654
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 18248 18970 18276 19790
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18524 18766 18552 19246
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18086 18552 18702
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18144 16584 18196 16590
rect 18064 16544 18144 16572
rect 18064 15502 18092 16544
rect 18144 16526 18196 16532
rect 18248 16266 18276 16594
rect 18420 16584 18472 16590
rect 18418 16552 18420 16561
rect 18472 16552 18474 16561
rect 18474 16510 18552 16538
rect 18418 16487 18474 16496
rect 18156 16238 18276 16266
rect 18156 16046 18184 16238
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15026 18092 15438
rect 18248 15162 18276 16118
rect 18524 15978 18552 16510
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18064 14618 18092 14962
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18432 14346 18460 14758
rect 18524 14550 18552 14826
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18420 14340 18472 14346
rect 18420 14282 18472 14288
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17512 12736 17632 12764
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17077 11996 17385 12005
rect 17077 11994 17083 11996
rect 17139 11994 17163 11996
rect 17219 11994 17243 11996
rect 17299 11994 17323 11996
rect 17379 11994 17385 11996
rect 17139 11942 17141 11994
rect 17321 11942 17323 11994
rect 17077 11940 17083 11942
rect 17139 11940 17163 11942
rect 17219 11940 17243 11942
rect 17299 11940 17323 11942
rect 17379 11940 17385 11942
rect 17077 11931 17385 11940
rect 17314 11112 17370 11121
rect 17314 11047 17316 11056
rect 17368 11047 17370 11056
rect 17316 11018 17368 11024
rect 17077 10908 17385 10917
rect 17077 10906 17083 10908
rect 17139 10906 17163 10908
rect 17219 10906 17243 10908
rect 17299 10906 17323 10908
rect 17379 10906 17385 10908
rect 17139 10854 17141 10906
rect 17321 10854 17323 10906
rect 17077 10852 17083 10854
rect 17139 10852 17163 10854
rect 17219 10852 17243 10854
rect 17299 10852 17323 10854
rect 17379 10852 17385 10854
rect 17077 10843 17385 10852
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17236 10606 17264 10678
rect 17224 10600 17276 10606
rect 17130 10568 17186 10577
rect 17224 10542 17276 10548
rect 17130 10503 17186 10512
rect 17144 10266 17172 10503
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17236 9926 17264 10542
rect 17420 10010 17448 12242
rect 17512 11642 17540 12736
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 11762 17632 12582
rect 17696 12306 17724 13466
rect 17880 13394 17908 13670
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12850 17908 13330
rect 17972 12986 18000 13874
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 18064 12714 18092 13262
rect 18432 13190 18460 14282
rect 18524 13190 18552 14486
rect 18616 13530 18644 20198
rect 18892 19990 18920 20295
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18786 19272 18842 19281
rect 18786 19207 18842 19216
rect 18800 18834 18828 19207
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18984 18057 19012 21830
rect 19352 21146 19380 22066
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19536 21690 19564 21898
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 19922 19380 20810
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19340 19440 19392 19446
rect 19444 19417 19472 21422
rect 19812 20398 19840 23666
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19340 19382 19392 19388
rect 19430 19408 19486 19417
rect 19352 18970 19380 19382
rect 19430 19343 19486 19352
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 18850 19472 19110
rect 19352 18834 19472 18850
rect 19628 18834 19656 19654
rect 19812 19514 19840 19654
rect 19904 19514 19932 24568
rect 20088 24342 20116 25366
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 21008 24954 21036 25162
rect 20996 24948 21048 24954
rect 20996 24890 21048 24896
rect 21192 24886 21220 25638
rect 21468 25226 21496 25638
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 21180 24880 21232 24886
rect 21086 24848 21142 24857
rect 21180 24822 21232 24828
rect 21086 24783 21142 24792
rect 21364 24812 21416 24818
rect 21100 24750 21128 24783
rect 21364 24754 21416 24760
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 21376 24410 21404 24754
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19996 23730 20024 24142
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19996 23186 20024 23666
rect 20088 23254 20116 24278
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21376 23866 21404 24142
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21468 23866 21496 24006
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 20732 23322 20760 23666
rect 20904 23656 20956 23662
rect 21284 23633 21312 23666
rect 21560 23662 21588 25706
rect 21548 23656 21600 23662
rect 20904 23598 20956 23604
rect 21270 23624 21326 23633
rect 20916 23322 20944 23598
rect 21548 23598 21600 23604
rect 21270 23559 21326 23568
rect 21560 23526 21588 23598
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19996 21962 20024 22374
rect 20548 22094 20576 23054
rect 20640 22166 20668 23122
rect 21008 22710 21036 23462
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20732 22234 20760 22510
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20628 22160 20680 22166
rect 20628 22102 20680 22108
rect 20456 22066 20576 22094
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19800 19508 19852 19514
rect 19800 19450 19852 19456
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19904 19394 19932 19450
rect 19812 19366 19932 19394
rect 19340 18828 19472 18834
rect 19392 18822 19472 18828
rect 19616 18828 19668 18834
rect 19340 18770 19392 18776
rect 19616 18770 19668 18776
rect 19352 18290 19380 18770
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 18970 18048 19026 18057
rect 18970 17983 19026 17992
rect 19444 17882 19472 18702
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19628 17542 19656 17818
rect 19812 17610 19840 19366
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19904 18970 19932 19246
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19904 17746 19932 18634
rect 19996 18426 20024 18906
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18708 16658 18736 16934
rect 18970 16688 19026 16697
rect 18696 16652 18748 16658
rect 18970 16623 19026 16632
rect 18696 16594 18748 16600
rect 18708 14958 18736 16594
rect 18984 16250 19012 16623
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15434 18828 15982
rect 19076 15706 19104 16390
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18892 15366 18920 15574
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 19168 15162 19196 17138
rect 19628 17105 19656 17478
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19614 17096 19670 17105
rect 19614 17031 19670 17040
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19352 15910 19380 16050
rect 19444 15910 19472 16458
rect 19628 16114 19656 16934
rect 19812 16794 19840 17138
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19812 16114 19840 16526
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 19352 14906 19380 15846
rect 19444 15026 19472 15846
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19628 14958 19656 15914
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15706 19932 15846
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19812 15162 19840 15370
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19524 14952 19576 14958
rect 19352 14900 19524 14906
rect 19352 14894 19576 14900
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19352 14878 19564 14894
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 13870 19748 14350
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18340 12442 18368 12718
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18432 12322 18460 13126
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 18340 12294 18460 12322
rect 17684 12096 17736 12102
rect 17868 12096 17920 12102
rect 17736 12056 17816 12084
rect 17684 12038 17736 12044
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17512 11614 17632 11642
rect 17420 9982 17540 10010
rect 17224 9920 17276 9926
rect 16946 9888 17002 9897
rect 17224 9862 17276 9868
rect 16946 9823 17002 9832
rect 17077 9820 17385 9829
rect 17077 9818 17083 9820
rect 17139 9818 17163 9820
rect 17219 9818 17243 9820
rect 17299 9818 17323 9820
rect 17379 9818 17385 9820
rect 17139 9766 17141 9818
rect 17321 9766 17323 9818
rect 17077 9764 17083 9766
rect 17139 9764 17163 9766
rect 17219 9764 17243 9766
rect 17299 9764 17323 9766
rect 17379 9764 17385 9766
rect 17077 9755 17385 9764
rect 17512 9722 17540 9982
rect 17500 9716 17552 9722
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16684 9450 16712 9687
rect 16776 9676 16988 9704
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16417 9276 16725 9285
rect 16417 9274 16423 9276
rect 16479 9274 16503 9276
rect 16559 9274 16583 9276
rect 16639 9274 16663 9276
rect 16719 9274 16725 9276
rect 16479 9222 16481 9274
rect 16661 9222 16663 9274
rect 16417 9220 16423 9222
rect 16479 9220 16503 9222
rect 16559 9220 16583 9222
rect 16639 9220 16663 9222
rect 16719 9220 16725 9222
rect 16417 9211 16725 9220
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8514 16712 8910
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8634 16804 8774
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16684 8486 16804 8514
rect 16417 8188 16725 8197
rect 16417 8186 16423 8188
rect 16479 8186 16503 8188
rect 16559 8186 16583 8188
rect 16639 8186 16663 8188
rect 16719 8186 16725 8188
rect 16479 8134 16481 8186
rect 16661 8134 16663 8186
rect 16417 8132 16423 8134
rect 16479 8132 16503 8134
rect 16559 8132 16583 8134
rect 16639 8132 16663 8134
rect 16719 8132 16725 8134
rect 16417 8123 16725 8132
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 7546 16620 7822
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 15752 6248 15804 6254
rect 15672 6208 15752 6236
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15580 5710 15608 6122
rect 15672 5846 15700 6208
rect 15752 6190 15804 6196
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15488 5324 15608 5352
rect 15476 5234 15528 5240
rect 15476 5176 15528 5182
rect 15488 5148 15516 5176
rect 15580 5166 15608 5324
rect 15396 5120 15516 5148
rect 15568 5160 15620 5166
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4758 14964 4966
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15396 4622 15424 5120
rect 15568 5102 15620 5108
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 15304 4146 15332 4558
rect 15488 4554 15516 4966
rect 15580 4729 15608 5102
rect 15566 4720 15622 4729
rect 15566 4655 15622 4664
rect 15672 4622 15700 5510
rect 15764 4826 15792 5714
rect 15856 5710 15884 6394
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15764 4690 15792 4762
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14292 3194 14320 3878
rect 15028 3602 15056 4014
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13912 2576 13964 2582
rect 13740 2524 13912 2530
rect 13740 2518 13964 2524
rect 13740 2502 13952 2518
rect 14568 2446 14596 3470
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3126 14964 3334
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15120 2650 15148 3470
rect 15580 3194 15608 4558
rect 15672 4010 15700 4558
rect 15856 4486 15884 5646
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15198 2680 15254 2689
rect 15108 2644 15160 2650
rect 15198 2615 15254 2624
rect 15108 2586 15160 2592
rect 15212 2446 15240 2615
rect 15396 2446 15424 2790
rect 15488 2446 15516 2926
rect 13820 2440 13872 2446
rect 13556 2400 13820 2428
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13556 800 13584 2400
rect 13820 2382 13872 2388
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15672 2378 15700 3606
rect 15948 2514 15976 7278
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6322 16160 6598
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16224 5710 16252 6734
rect 16316 6730 16344 7142
rect 16417 7100 16725 7109
rect 16417 7098 16423 7100
rect 16479 7098 16503 7100
rect 16559 7098 16583 7100
rect 16639 7098 16663 7100
rect 16719 7098 16725 7100
rect 16479 7046 16481 7098
rect 16661 7046 16663 7098
rect 16417 7044 16423 7046
rect 16479 7044 16503 7046
rect 16559 7044 16583 7046
rect 16639 7044 16663 7046
rect 16719 7044 16725 7046
rect 16417 7035 16725 7044
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16316 6458 16344 6666
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 5704 16264 5710
rect 16316 5681 16344 6258
rect 16408 6118 16436 6394
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16417 6012 16725 6021
rect 16417 6010 16423 6012
rect 16479 6010 16503 6012
rect 16559 6010 16583 6012
rect 16639 6010 16663 6012
rect 16719 6010 16725 6012
rect 16479 5958 16481 6010
rect 16661 5958 16663 6010
rect 16417 5956 16423 5958
rect 16479 5956 16503 5958
rect 16559 5956 16583 5958
rect 16639 5956 16663 5958
rect 16719 5956 16725 5958
rect 16417 5947 16725 5956
rect 16212 5646 16264 5652
rect 16302 5672 16358 5681
rect 16302 5607 16358 5616
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16026 5264 16082 5273
rect 16500 5234 16528 5510
rect 16776 5370 16804 8486
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16026 5199 16028 5208
rect 16080 5199 16082 5208
rect 16488 5228 16540 5234
rect 16028 5170 16080 5176
rect 16488 5170 16540 5176
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16040 4826 16068 4966
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16132 3466 16160 4966
rect 16316 4826 16344 4966
rect 16417 4924 16725 4933
rect 16417 4922 16423 4924
rect 16479 4922 16503 4924
rect 16559 4922 16583 4924
rect 16639 4922 16663 4924
rect 16719 4922 16725 4924
rect 16479 4870 16481 4922
rect 16661 4870 16663 4922
rect 16417 4868 16423 4870
rect 16479 4868 16503 4870
rect 16559 4868 16583 4870
rect 16639 4868 16663 4870
rect 16719 4868 16725 4870
rect 16417 4859 16725 4868
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16396 4752 16448 4758
rect 16394 4720 16396 4729
rect 16448 4720 16450 4729
rect 16394 4655 16450 4664
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16417 3836 16725 3845
rect 16417 3834 16423 3836
rect 16479 3834 16503 3836
rect 16559 3834 16583 3836
rect 16639 3834 16663 3836
rect 16719 3834 16725 3836
rect 16479 3782 16481 3834
rect 16661 3782 16663 3834
rect 16417 3780 16423 3782
rect 16479 3780 16503 3782
rect 16559 3780 16583 3782
rect 16639 3780 16663 3782
rect 16719 3780 16725 3782
rect 16417 3771 16725 3780
rect 16776 3602 16804 4558
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16868 2854 16896 9046
rect 16960 7546 16988 9676
rect 17038 9688 17094 9697
rect 17500 9658 17552 9664
rect 17038 9623 17094 9632
rect 17052 9450 17080 9623
rect 17604 9602 17632 11614
rect 17788 9897 17816 12056
rect 17868 12038 17920 12044
rect 17880 11218 17908 12038
rect 18340 11830 18368 12294
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11286 18000 11494
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17774 9888 17830 9897
rect 17774 9823 17830 9832
rect 17682 9688 17738 9697
rect 17972 9674 18000 11222
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18064 9722 18092 10746
rect 17682 9623 17738 9632
rect 17926 9646 18000 9674
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17512 9574 17632 9602
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 17052 8974 17080 9386
rect 17512 9058 17540 9574
rect 17696 9110 17724 9623
rect 17926 9602 17954 9646
rect 17788 9574 17954 9602
rect 18236 9580 18288 9586
rect 17684 9104 17736 9110
rect 17512 9030 17632 9058
rect 17684 9046 17736 9052
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17077 8732 17385 8741
rect 17077 8730 17083 8732
rect 17139 8730 17163 8732
rect 17219 8730 17243 8732
rect 17299 8730 17323 8732
rect 17379 8730 17385 8732
rect 17139 8678 17141 8730
rect 17321 8678 17323 8730
rect 17077 8676 17083 8678
rect 17139 8676 17163 8678
rect 17219 8676 17243 8678
rect 17299 8676 17323 8678
rect 17379 8676 17385 8678
rect 17077 8667 17385 8676
rect 17512 8430 17540 8774
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17236 7954 17264 8366
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17077 7644 17385 7653
rect 17077 7642 17083 7644
rect 17139 7642 17163 7644
rect 17219 7642 17243 7644
rect 17299 7642 17323 7644
rect 17379 7642 17385 7644
rect 17139 7590 17141 7642
rect 17321 7590 17323 7642
rect 17077 7588 17083 7590
rect 17139 7588 17163 7590
rect 17219 7588 17243 7590
rect 17299 7588 17323 7590
rect 17379 7588 17385 7590
rect 17077 7579 17385 7588
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 5914 16988 6734
rect 17077 6556 17385 6565
rect 17077 6554 17083 6556
rect 17139 6554 17163 6556
rect 17219 6554 17243 6556
rect 17299 6554 17323 6556
rect 17379 6554 17385 6556
rect 17139 6502 17141 6554
rect 17321 6502 17323 6554
rect 17077 6500 17083 6502
rect 17139 6500 17163 6502
rect 17219 6500 17243 6502
rect 17299 6500 17323 6502
rect 17379 6500 17385 6502
rect 17077 6491 17385 6500
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17144 5846 17172 6054
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17236 5710 17264 5850
rect 17328 5710 17356 6190
rect 17132 5704 17184 5710
rect 17130 5672 17132 5681
rect 17224 5704 17276 5710
rect 17184 5672 17186 5681
rect 17224 5646 17276 5652
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17130 5607 17186 5616
rect 17077 5468 17385 5477
rect 17077 5466 17083 5468
rect 17139 5466 17163 5468
rect 17219 5466 17243 5468
rect 17299 5466 17323 5468
rect 17379 5466 17385 5468
rect 17139 5414 17141 5466
rect 17321 5414 17323 5466
rect 17077 5412 17083 5414
rect 17139 5412 17163 5414
rect 17219 5412 17243 5414
rect 17299 5412 17323 5414
rect 17379 5412 17385 5414
rect 17077 5403 17385 5412
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16417 2748 16725 2757
rect 16417 2746 16423 2748
rect 16479 2746 16503 2748
rect 16559 2746 16583 2748
rect 16639 2746 16663 2748
rect 16719 2746 16725 2748
rect 16479 2694 16481 2746
rect 16661 2694 16663 2746
rect 16417 2692 16423 2694
rect 16479 2692 16503 2694
rect 16559 2692 16583 2694
rect 16639 2692 16663 2694
rect 16719 2692 16725 2694
rect 16417 2683 16725 2692
rect 16960 2666 16988 5306
rect 17420 5302 17448 7210
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17077 4380 17385 4389
rect 17077 4378 17083 4380
rect 17139 4378 17163 4380
rect 17219 4378 17243 4380
rect 17299 4378 17323 4380
rect 17379 4378 17385 4380
rect 17139 4326 17141 4378
rect 17321 4326 17323 4378
rect 17077 4324 17083 4326
rect 17139 4324 17163 4326
rect 17219 4324 17243 4326
rect 17299 4324 17323 4326
rect 17379 4324 17385 4326
rect 17077 4315 17385 4324
rect 17512 4010 17540 7958
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17077 3292 17385 3301
rect 17077 3290 17083 3292
rect 17139 3290 17163 3292
rect 17219 3290 17243 3292
rect 17299 3290 17323 3292
rect 17379 3290 17385 3292
rect 17139 3238 17141 3290
rect 17321 3238 17323 3290
rect 17077 3236 17083 3238
rect 17139 3236 17163 3238
rect 17219 3236 17243 3238
rect 17299 3236 17323 3238
rect 17379 3236 17385 3238
rect 17077 3227 17385 3236
rect 17420 3194 17448 3402
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17512 2922 17540 3946
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 16776 2638 16988 2666
rect 17052 2650 17080 2858
rect 17040 2644 17092 2650
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16776 2446 16804 2638
rect 17040 2586 17092 2592
rect 17604 2496 17632 9030
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 8634 17724 8910
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17788 8022 17816 9574
rect 18236 9522 18288 9528
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 8090 18000 8910
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8566 18092 8774
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7313 17724 7686
rect 17682 7304 17738 7313
rect 17682 7239 17738 7248
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17696 6186 17724 7142
rect 17788 6798 17816 7754
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17774 6624 17830 6633
rect 17774 6559 17830 6568
rect 17684 6180 17736 6186
rect 17684 6122 17736 6128
rect 17788 6066 17816 6559
rect 17696 6038 17816 6066
rect 17880 6168 17908 7822
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17972 6934 18000 7482
rect 18064 7410 18092 8230
rect 18156 8090 18184 8570
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18064 6798 18092 6938
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18156 6644 18184 7346
rect 17972 6616 18184 6644
rect 17972 6361 18000 6616
rect 18052 6384 18104 6390
rect 17958 6352 18014 6361
rect 18052 6326 18104 6332
rect 17958 6287 18014 6296
rect 17960 6180 18012 6186
rect 17880 6140 17960 6168
rect 17696 4146 17724 6038
rect 17880 5370 17908 6140
rect 17960 6122 18012 6128
rect 18064 5710 18092 6326
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17880 4690 17908 5306
rect 18248 5302 18276 9522
rect 18340 9466 18368 11766
rect 18524 11626 18552 13126
rect 18616 12918 18644 13466
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18616 12306 18644 12854
rect 18892 12782 18920 13194
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12918 19380 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18892 12374 18920 12718
rect 19444 12442 19472 13262
rect 19812 12782 19840 14894
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10062 18460 10950
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18340 9438 18460 9466
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18340 7342 18368 9318
rect 18432 8090 18460 9438
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18340 6390 18368 7142
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18432 6254 18460 7754
rect 18524 7546 18552 11562
rect 18708 11150 18736 12242
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18800 11150 18828 11562
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18708 10810 18736 11086
rect 18892 10810 18920 11290
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19614 10160 19670 10169
rect 19614 10095 19670 10104
rect 19628 10062 19656 10095
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 18800 9518 18828 9862
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18708 8430 18736 8978
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 7954 18736 8366
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18524 7002 18552 7346
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 18800 5234 18828 9454
rect 19260 8974 19288 9862
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18984 7002 19012 7346
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 4282 18000 4490
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 3126 17724 4082
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17788 2582 17816 3470
rect 18984 2582 19012 6734
rect 19260 6730 19288 7686
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19260 4826 19288 6666
rect 19352 6390 19380 7142
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5370 19564 5646
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19536 4146 19564 5306
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19536 3602 19564 4082
rect 19720 4078 19748 9862
rect 19812 9654 19840 10542
rect 19904 10266 19932 14826
rect 19996 14618 20024 14962
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13530 20024 13806
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 12850 20116 20198
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19812 9042 19840 9590
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19904 8634 19932 10202
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19904 7410 19932 8570
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19812 6458 19840 6802
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19812 5914 19840 6394
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 20088 5642 20116 6598
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19720 2774 19748 4014
rect 20180 2774 20208 21490
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20272 15094 20300 21354
rect 20456 20466 20484 22066
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21486 20576 21830
rect 20640 21486 20668 22102
rect 21284 22094 21312 22918
rect 21284 22066 21404 22094
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21284 21690 21312 21966
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20628 21072 20680 21078
rect 20628 21014 20680 21020
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 17490 20484 20402
rect 20548 19174 20576 20878
rect 20640 19990 20668 21014
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21192 20602 21220 20810
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18834 20576 19110
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20548 18290 20576 18770
rect 21008 18426 21036 19654
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21192 18698 21220 19178
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 17678 20576 18226
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 21284 17610 21312 18022
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 20456 17462 20576 17490
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20364 16590 20392 17138
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20364 16250 20392 16526
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20272 13394 20300 15030
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20456 12918 20484 14350
rect 20548 14278 20576 17462
rect 20824 17338 20852 17546
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 21376 17218 21404 22066
rect 21640 21548 21692 21554
rect 21640 21490 21692 21496
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21468 20874 21496 21286
rect 21652 21146 21680 21490
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 21456 20868 21508 20874
rect 21456 20810 21508 20816
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21560 18698 21588 19654
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21652 18426 21680 19314
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 21546 18048 21602 18057
rect 21546 17983 21602 17992
rect 21376 17190 21496 17218
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20640 16658 20668 17002
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16794 20944 16934
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 21192 16454 21220 17070
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15162 20760 15846
rect 20916 15706 20944 16390
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14482 20760 14758
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21008 13530 21036 13942
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20534 13288 20590 13297
rect 20534 13223 20536 13232
rect 20588 13223 20590 13232
rect 20536 13194 20588 13200
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 19444 2746 19748 2774
rect 20088 2746 20208 2774
rect 20272 2774 20300 12786
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20364 12442 20392 12718
rect 20352 12436 20404 12442
rect 20456 12434 20484 12854
rect 20456 12406 20576 12434
rect 20352 12378 20404 12384
rect 20364 11830 20392 12378
rect 20548 12306 20576 12406
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20456 11898 20484 12174
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20364 10130 20392 11766
rect 20640 11234 20668 13330
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 11626 20852 12650
rect 21100 12434 21128 15982
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21376 13530 21404 14282
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12986 21220 13262
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21008 12406 21128 12434
rect 21468 12434 21496 17190
rect 21560 14074 21588 17983
rect 21652 17134 21680 18090
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21560 12986 21588 13262
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21468 12406 21588 12434
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20548 11218 20668 11234
rect 20536 11212 20668 11218
rect 20588 11206 20668 11212
rect 20536 11154 20588 11160
rect 20824 11098 20852 11562
rect 20640 11070 20852 11098
rect 20640 10198 20668 11070
rect 20718 10704 20774 10713
rect 20718 10639 20774 10648
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 8566 20392 10066
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20364 6322 20392 8502
rect 20640 8362 20668 10134
rect 20732 10062 20760 10639
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 8634 20852 9522
rect 20916 9178 20944 9862
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20640 6984 20668 8298
rect 20732 7886 20760 8366
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20456 6956 20668 6984
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20364 5778 20392 6258
rect 20456 6186 20484 6956
rect 20732 6882 20760 7822
rect 21008 7546 21036 12406
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21468 11898 21496 12106
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21180 11144 21232 11150
rect 21376 11132 21404 11494
rect 21232 11104 21404 11132
rect 21180 11086 21232 11092
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10810 21128 10950
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20548 6854 20760 6882
rect 20548 6798 20576 6854
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20456 5846 20484 6122
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20364 5302 20392 5714
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20364 5166 20392 5238
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20456 5098 20484 5782
rect 20548 5710 20576 6734
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 5846 20760 6598
rect 20824 6458 20852 6666
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20824 5370 20852 6258
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20640 4826 20668 4966
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 20916 4214 20944 4422
rect 20904 4208 20956 4214
rect 20904 4150 20956 4156
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20916 3194 20944 3470
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21008 2990 21036 7482
rect 21100 5658 21128 10406
rect 21376 10130 21404 11104
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21192 9178 21220 9930
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21284 8974 21312 9318
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21284 7970 21312 8774
rect 21192 7954 21312 7970
rect 21180 7948 21312 7954
rect 21232 7942 21312 7948
rect 21180 7890 21232 7896
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21192 5778 21220 7142
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 21100 5630 21220 5658
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21100 4593 21128 5170
rect 21086 4584 21142 4593
rect 21086 4519 21142 4528
rect 21086 3088 21142 3097
rect 21192 3074 21220 5630
rect 21376 5166 21404 10066
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21468 6458 21496 6666
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21560 3398 21588 12406
rect 21652 9994 21680 14962
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21744 6662 21772 26250
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21836 21554 21864 23462
rect 21928 23186 21956 26250
rect 22848 25684 22876 26454
rect 22940 25906 22968 28591
rect 23202 28381 23258 29181
rect 23846 28506 23902 29181
rect 24490 28506 24546 29181
rect 23846 28478 23980 28506
rect 23846 28381 23902 28478
rect 23216 26586 23244 28381
rect 23952 26586 23980 28478
rect 24490 28478 24624 28506
rect 24490 28381 24546 28478
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 24596 26450 24624 28478
rect 25778 28381 25834 29181
rect 26422 28381 26478 29181
rect 25502 27976 25558 27985
rect 25502 27911 25558 27920
rect 24858 26616 24914 26625
rect 24858 26551 24914 26560
rect 24872 26518 24900 26551
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 23848 26308 23900 26314
rect 23848 26250 23900 26256
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23032 26042 23060 26182
rect 23020 26036 23072 26042
rect 23020 25978 23072 25984
rect 22928 25900 22980 25906
rect 22928 25842 22980 25848
rect 22848 25656 22968 25684
rect 22604 25596 22912 25605
rect 22604 25594 22610 25596
rect 22666 25594 22690 25596
rect 22746 25594 22770 25596
rect 22826 25594 22850 25596
rect 22906 25594 22912 25596
rect 22666 25542 22668 25594
rect 22848 25542 22850 25594
rect 22604 25540 22610 25542
rect 22666 25540 22690 25542
rect 22746 25540 22770 25542
rect 22826 25540 22850 25542
rect 22906 25540 22912 25542
rect 22604 25531 22912 25540
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 22020 23798 22048 24074
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22204 23662 22232 25094
rect 22604 24508 22912 24517
rect 22604 24506 22610 24508
rect 22666 24506 22690 24508
rect 22746 24506 22770 24508
rect 22826 24506 22850 24508
rect 22906 24506 22912 24508
rect 22666 24454 22668 24506
rect 22848 24454 22850 24506
rect 22604 24452 22610 24454
rect 22666 24452 22690 24454
rect 22746 24452 22770 24454
rect 22826 24452 22850 24454
rect 22906 24452 22912 24454
rect 22604 24443 22912 24452
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22604 23420 22912 23429
rect 22604 23418 22610 23420
rect 22666 23418 22690 23420
rect 22746 23418 22770 23420
rect 22826 23418 22850 23420
rect 22906 23418 22912 23420
rect 22666 23366 22668 23418
rect 22848 23366 22850 23418
rect 22604 23364 22610 23366
rect 22666 23364 22690 23366
rect 22746 23364 22770 23366
rect 22826 23364 22850 23366
rect 22906 23364 22912 23366
rect 22604 23355 22912 23364
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 21928 22778 21956 23122
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22604 22332 22912 22341
rect 22604 22330 22610 22332
rect 22666 22330 22690 22332
rect 22746 22330 22770 22332
rect 22826 22330 22850 22332
rect 22906 22330 22912 22332
rect 22666 22278 22668 22330
rect 22848 22278 22850 22330
rect 22604 22276 22610 22278
rect 22666 22276 22690 22278
rect 22746 22276 22770 22278
rect 22826 22276 22850 22278
rect 22906 22276 22912 22278
rect 22604 22267 22912 22276
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 22604 21244 22912 21253
rect 22604 21242 22610 21244
rect 22666 21242 22690 21244
rect 22746 21242 22770 21244
rect 22826 21242 22850 21244
rect 22906 21242 22912 21244
rect 22666 21190 22668 21242
rect 22848 21190 22850 21242
rect 22604 21188 22610 21190
rect 22666 21188 22690 21190
rect 22746 21188 22770 21190
rect 22826 21188 22850 21190
rect 22906 21188 22912 21190
rect 22604 21179 22912 21188
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20602 22232 20742
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19446 22232 20198
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 18426 22324 18566
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22388 18222 22416 20334
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22388 17762 22416 18158
rect 22480 17882 22508 20402
rect 22604 20156 22912 20165
rect 22604 20154 22610 20156
rect 22666 20154 22690 20156
rect 22746 20154 22770 20156
rect 22826 20154 22850 20156
rect 22906 20154 22912 20156
rect 22666 20102 22668 20154
rect 22848 20102 22850 20154
rect 22604 20100 22610 20102
rect 22666 20100 22690 20102
rect 22746 20100 22770 20102
rect 22826 20100 22850 20102
rect 22906 20100 22912 20102
rect 22604 20091 22912 20100
rect 22604 19068 22912 19077
rect 22604 19066 22610 19068
rect 22666 19066 22690 19068
rect 22746 19066 22770 19068
rect 22826 19066 22850 19068
rect 22906 19066 22912 19068
rect 22666 19014 22668 19066
rect 22848 19014 22850 19066
rect 22604 19012 22610 19014
rect 22666 19012 22690 19014
rect 22746 19012 22770 19014
rect 22826 19012 22850 19014
rect 22906 19012 22912 19014
rect 22604 19003 22912 19012
rect 22604 17980 22912 17989
rect 22604 17978 22610 17980
rect 22666 17978 22690 17980
rect 22746 17978 22770 17980
rect 22826 17978 22850 17980
rect 22906 17978 22912 17980
rect 22666 17926 22668 17978
rect 22848 17926 22850 17978
rect 22604 17924 22610 17926
rect 22666 17924 22690 17926
rect 22746 17924 22770 17926
rect 22826 17924 22850 17926
rect 22906 17924 22912 17926
rect 22604 17915 22912 17924
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22204 17746 22416 17762
rect 22192 17740 22416 17746
rect 22244 17734 22416 17740
rect 22192 17682 22244 17688
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 16590 21864 17478
rect 22388 17134 22416 17734
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22664 17338 22692 17478
rect 22848 17338 22876 17546
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22604 16892 22912 16901
rect 22604 16890 22610 16892
rect 22666 16890 22690 16892
rect 22746 16890 22770 16892
rect 22826 16890 22850 16892
rect 22906 16890 22912 16892
rect 22666 16838 22668 16890
rect 22848 16838 22850 16890
rect 22604 16836 22610 16838
rect 22666 16836 22690 16838
rect 22746 16836 22770 16838
rect 22826 16836 22850 16838
rect 22906 16836 22912 16838
rect 22604 16827 22912 16836
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21836 16182 21864 16526
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21928 16114 21956 16730
rect 22192 16720 22244 16726
rect 22376 16720 22428 16726
rect 22192 16662 22244 16668
rect 22296 16680 22376 16708
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22020 16250 22048 16390
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22020 14890 22048 15302
rect 22112 14890 22140 15982
rect 22204 15978 22232 16662
rect 22296 16522 22324 16680
rect 22376 16662 22428 16668
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22374 16008 22430 16017
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22284 15972 22336 15978
rect 22374 15943 22430 15952
rect 22284 15914 22336 15920
rect 22204 15706 22232 15914
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 21916 14816 21968 14822
rect 22204 14770 22232 15642
rect 22296 15570 22324 15914
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22296 15434 22324 15506
rect 22284 15428 22336 15434
rect 22284 15370 22336 15376
rect 22296 15008 22324 15370
rect 22388 15162 22416 15943
rect 22480 15434 22508 16390
rect 22848 16250 22876 16458
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22604 15804 22912 15813
rect 22604 15802 22610 15804
rect 22666 15802 22690 15804
rect 22746 15802 22770 15804
rect 22826 15802 22850 15804
rect 22906 15802 22912 15804
rect 22666 15750 22668 15802
rect 22848 15750 22850 15802
rect 22604 15748 22610 15750
rect 22666 15748 22690 15750
rect 22746 15748 22770 15750
rect 22826 15748 22850 15750
rect 22906 15748 22912 15750
rect 22604 15739 22912 15748
rect 22468 15428 22520 15434
rect 22468 15370 22520 15376
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22376 15020 22428 15026
rect 22296 14980 22376 15008
rect 22376 14962 22428 14968
rect 22940 14906 22968 25656
rect 23124 20466 23152 26182
rect 23264 26140 23572 26149
rect 23264 26138 23270 26140
rect 23326 26138 23350 26140
rect 23406 26138 23430 26140
rect 23486 26138 23510 26140
rect 23566 26138 23572 26140
rect 23326 26086 23328 26138
rect 23508 26086 23510 26138
rect 23264 26084 23270 26086
rect 23326 26084 23350 26086
rect 23406 26084 23430 26086
rect 23486 26084 23510 26086
rect 23566 26084 23572 26086
rect 23264 26075 23572 26084
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23264 25052 23572 25061
rect 23264 25050 23270 25052
rect 23326 25050 23350 25052
rect 23406 25050 23430 25052
rect 23486 25050 23510 25052
rect 23566 25050 23572 25052
rect 23326 24998 23328 25050
rect 23508 24998 23510 25050
rect 23264 24996 23270 24998
rect 23326 24996 23350 24998
rect 23406 24996 23430 24998
rect 23486 24996 23510 24998
rect 23566 24996 23572 24998
rect 23264 24987 23572 24996
rect 23264 23964 23572 23973
rect 23264 23962 23270 23964
rect 23326 23962 23350 23964
rect 23406 23962 23430 23964
rect 23486 23962 23510 23964
rect 23566 23962 23572 23964
rect 23326 23910 23328 23962
rect 23508 23910 23510 23962
rect 23264 23908 23270 23910
rect 23326 23908 23350 23910
rect 23406 23908 23430 23910
rect 23486 23908 23510 23910
rect 23566 23908 23572 23910
rect 23264 23899 23572 23908
rect 23768 23526 23796 25094
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23264 22876 23572 22885
rect 23264 22874 23270 22876
rect 23326 22874 23350 22876
rect 23406 22874 23430 22876
rect 23486 22874 23510 22876
rect 23566 22874 23572 22876
rect 23326 22822 23328 22874
rect 23508 22822 23510 22874
rect 23264 22820 23270 22822
rect 23326 22820 23350 22822
rect 23406 22820 23430 22822
rect 23486 22820 23510 22822
rect 23566 22820 23572 22822
rect 23264 22811 23572 22820
rect 23860 22094 23888 26250
rect 25318 25936 25374 25945
rect 25318 25871 25320 25880
rect 25372 25871 25374 25880
rect 25320 25842 25372 25848
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23768 22066 23888 22094
rect 23264 21788 23572 21797
rect 23264 21786 23270 21788
rect 23326 21786 23350 21788
rect 23406 21786 23430 21788
rect 23486 21786 23510 21788
rect 23566 21786 23572 21788
rect 23326 21734 23328 21786
rect 23508 21734 23510 21786
rect 23264 21732 23270 21734
rect 23326 21732 23350 21734
rect 23406 21732 23430 21734
rect 23486 21732 23510 21734
rect 23566 21732 23572 21734
rect 23264 21723 23572 21732
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23264 20700 23572 20709
rect 23264 20698 23270 20700
rect 23326 20698 23350 20700
rect 23406 20698 23430 20700
rect 23486 20698 23510 20700
rect 23566 20698 23572 20700
rect 23326 20646 23328 20698
rect 23508 20646 23510 20698
rect 23264 20644 23270 20646
rect 23326 20644 23350 20646
rect 23406 20644 23430 20646
rect 23486 20644 23510 20646
rect 23566 20644 23572 20646
rect 23264 20635 23572 20644
rect 23676 20602 23704 21286
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23124 19514 23152 19654
rect 23264 19612 23572 19621
rect 23264 19610 23270 19612
rect 23326 19610 23350 19612
rect 23406 19610 23430 19612
rect 23486 19610 23510 19612
rect 23566 19610 23572 19612
rect 23326 19558 23328 19610
rect 23508 19558 23510 19610
rect 23264 19556 23270 19558
rect 23326 19556 23350 19558
rect 23406 19556 23430 19558
rect 23486 19556 23510 19558
rect 23566 19556 23572 19558
rect 23264 19547 23572 19556
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 23676 19446 23704 20198
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23032 18766 23060 19246
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 23032 18222 23060 18702
rect 23124 18426 23152 19110
rect 23492 18834 23520 19178
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23264 18524 23572 18533
rect 23264 18522 23270 18524
rect 23326 18522 23350 18524
rect 23406 18522 23430 18524
rect 23486 18522 23510 18524
rect 23566 18522 23572 18524
rect 23326 18470 23328 18522
rect 23508 18470 23510 18522
rect 23264 18468 23270 18470
rect 23326 18468 23350 18470
rect 23406 18468 23430 18470
rect 23486 18468 23510 18470
rect 23566 18468 23572 18470
rect 23264 18459 23572 18468
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23032 15978 23060 18158
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23216 17524 23244 17818
rect 23308 17678 23336 18294
rect 23676 17746 23704 18770
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23124 17496 23244 17524
rect 23124 17338 23152 17496
rect 23264 17436 23572 17445
rect 23264 17434 23270 17436
rect 23326 17434 23350 17436
rect 23406 17434 23430 17436
rect 23486 17434 23510 17436
rect 23566 17434 23572 17436
rect 23326 17382 23328 17434
rect 23508 17382 23510 17434
rect 23264 17380 23270 17382
rect 23326 17380 23350 17382
rect 23406 17380 23430 17382
rect 23486 17380 23510 17382
rect 23566 17380 23572 17382
rect 23264 17371 23572 17380
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23676 17270 23704 17682
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23676 16726 23704 17206
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23264 16348 23572 16357
rect 23264 16346 23270 16348
rect 23326 16346 23350 16348
rect 23406 16346 23430 16348
rect 23486 16346 23510 16348
rect 23566 16346 23572 16348
rect 23326 16294 23328 16346
rect 23508 16294 23510 16346
rect 23264 16292 23270 16294
rect 23326 16292 23350 16294
rect 23406 16292 23430 16294
rect 23486 16292 23510 16294
rect 23566 16292 23572 16294
rect 23264 16283 23572 16292
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23400 16153 23428 16186
rect 23202 16144 23258 16153
rect 23202 16079 23204 16088
rect 23256 16079 23258 16088
rect 23386 16144 23442 16153
rect 23768 16130 23796 22066
rect 23846 19816 23902 19825
rect 23846 19751 23848 19760
rect 23900 19751 23902 19760
rect 23848 19722 23900 19728
rect 23952 18986 23980 25638
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24492 25288 24544 25294
rect 24872 25265 24900 25434
rect 24492 25230 24544 25236
rect 24858 25256 24914 25265
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23860 18958 23980 18986
rect 23860 16658 23888 18958
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 23952 17814 23980 18838
rect 23940 17808 23992 17814
rect 23940 17750 23992 17756
rect 23952 17066 23980 17750
rect 24044 17678 24072 25094
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24136 19922 24164 21422
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23860 16250 23888 16390
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23768 16102 23888 16130
rect 23386 16079 23442 16088
rect 23204 16050 23256 16056
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23020 15972 23072 15978
rect 23020 15914 23072 15920
rect 23400 15706 23428 15982
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23264 15260 23572 15269
rect 23264 15258 23270 15260
rect 23326 15258 23350 15260
rect 23406 15258 23430 15260
rect 23486 15258 23510 15260
rect 23566 15258 23572 15260
rect 23326 15206 23328 15258
rect 23508 15206 23510 15258
rect 23264 15204 23270 15206
rect 23326 15204 23350 15206
rect 23406 15204 23430 15206
rect 23486 15204 23510 15206
rect 23566 15204 23572 15206
rect 23264 15195 23572 15204
rect 23388 14952 23440 14958
rect 22376 14884 22428 14890
rect 22940 14878 23060 14906
rect 23388 14894 23440 14900
rect 22376 14826 22428 14832
rect 21916 14758 21968 14764
rect 21928 14618 21956 14758
rect 22020 14742 22232 14770
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12434 21956 13126
rect 21836 12406 21956 12434
rect 21836 10010 21864 12406
rect 21928 12374 21956 12406
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10198 21956 11018
rect 22020 10962 22048 14742
rect 22190 14376 22246 14385
rect 22190 14311 22246 14320
rect 22204 14278 22232 14311
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22112 11082 22140 12106
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22020 10934 22140 10962
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22020 10266 22048 10610
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21836 9982 21956 10010
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21744 5914 21772 6258
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21836 5642 21864 6054
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21142 3046 21220 3074
rect 21744 3058 21772 5102
rect 21272 3052 21324 3058
rect 21086 3023 21142 3032
rect 21272 2994 21324 3000
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 20272 2746 20484 2774
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 17684 2508 17736 2514
rect 17604 2468 17684 2496
rect 17684 2450 17736 2456
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16856 2440 16908 2446
rect 19444 2417 19472 2746
rect 20088 2666 20116 2746
rect 20088 2638 20392 2666
rect 20364 2582 20392 2638
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 20456 2446 20484 2746
rect 21284 2650 21312 2994
rect 21928 2774 21956 9982
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22020 8362 22048 8774
rect 22112 8378 22140 10934
rect 22204 9874 22232 14214
rect 22388 11898 22416 14826
rect 22604 14716 22912 14725
rect 22604 14714 22610 14716
rect 22666 14714 22690 14716
rect 22746 14714 22770 14716
rect 22826 14714 22850 14716
rect 22906 14714 22912 14716
rect 22666 14662 22668 14714
rect 22848 14662 22850 14714
rect 22604 14660 22610 14662
rect 22666 14660 22690 14662
rect 22746 14660 22770 14662
rect 22826 14660 22850 14662
rect 22906 14660 22912 14662
rect 22604 14651 22912 14660
rect 22604 13628 22912 13637
rect 22604 13626 22610 13628
rect 22666 13626 22690 13628
rect 22746 13626 22770 13628
rect 22826 13626 22850 13628
rect 22906 13626 22912 13628
rect 22666 13574 22668 13626
rect 22848 13574 22850 13626
rect 22604 13572 22610 13574
rect 22666 13572 22690 13574
rect 22746 13572 22770 13574
rect 22826 13572 22850 13574
rect 22906 13572 22912 13574
rect 22604 13563 22912 13572
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22604 12540 22912 12549
rect 22604 12538 22610 12540
rect 22666 12538 22690 12540
rect 22746 12538 22770 12540
rect 22826 12538 22850 12540
rect 22906 12538 22912 12540
rect 22666 12486 22668 12538
rect 22848 12486 22850 12538
rect 22604 12484 22610 12486
rect 22666 12484 22690 12486
rect 22746 12484 22770 12486
rect 22826 12484 22850 12486
rect 22906 12484 22912 12486
rect 22604 12475 22912 12484
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 10470 22324 11630
rect 22604 11452 22912 11461
rect 22604 11450 22610 11452
rect 22666 11450 22690 11452
rect 22746 11450 22770 11452
rect 22826 11450 22850 11452
rect 22906 11450 22912 11452
rect 22666 11398 22668 11450
rect 22848 11398 22850 11450
rect 22604 11396 22610 11398
rect 22666 11396 22690 11398
rect 22746 11396 22770 11398
rect 22826 11396 22850 11398
rect 22906 11396 22912 11398
rect 22604 11387 22912 11396
rect 22940 11354 22968 12718
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23032 11234 23060 14878
rect 23400 14618 23428 14894
rect 23768 14618 23796 15506
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23264 14172 23572 14181
rect 23264 14170 23270 14172
rect 23326 14170 23350 14172
rect 23406 14170 23430 14172
rect 23486 14170 23510 14172
rect 23566 14170 23572 14172
rect 23326 14118 23328 14170
rect 23508 14118 23510 14170
rect 23264 14116 23270 14118
rect 23326 14116 23350 14118
rect 23406 14116 23430 14118
rect 23486 14116 23510 14118
rect 23566 14116 23572 14118
rect 23264 14107 23572 14116
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23264 13084 23572 13093
rect 23264 13082 23270 13084
rect 23326 13082 23350 13084
rect 23406 13082 23430 13084
rect 23486 13082 23510 13084
rect 23566 13082 23572 13084
rect 23326 13030 23328 13082
rect 23508 13030 23510 13082
rect 23264 13028 23270 13030
rect 23326 13028 23350 13030
rect 23406 13028 23430 13030
rect 23486 13028 23510 13030
rect 23566 13028 23572 13030
rect 23264 13019 23572 13028
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 22940 11206 23060 11234
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22604 10364 22912 10373
rect 22604 10362 22610 10364
rect 22666 10362 22690 10364
rect 22746 10362 22770 10364
rect 22826 10362 22850 10364
rect 22906 10362 22912 10364
rect 22666 10310 22668 10362
rect 22848 10310 22850 10362
rect 22604 10308 22610 10310
rect 22666 10308 22690 10310
rect 22746 10308 22770 10310
rect 22826 10308 22850 10310
rect 22906 10308 22912 10310
rect 22604 10299 22912 10308
rect 22744 10260 22796 10266
rect 22940 10248 22968 11206
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23032 10266 23060 11086
rect 23124 10674 23152 12922
rect 23676 12918 23704 13126
rect 23768 12986 23796 13806
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23860 12306 23888 16102
rect 23952 15706 23980 16526
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 15473 23980 15506
rect 23938 15464 23994 15473
rect 23938 15399 23994 15408
rect 24044 14006 24072 16934
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23952 12442 23980 13262
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 24032 12368 24084 12374
rect 24032 12310 24084 12316
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23264 11996 23572 12005
rect 23264 11994 23270 11996
rect 23326 11994 23350 11996
rect 23406 11994 23430 11996
rect 23486 11994 23510 11996
rect 23566 11994 23572 11996
rect 23326 11942 23328 11994
rect 23508 11942 23510 11994
rect 23264 11940 23270 11942
rect 23326 11940 23350 11942
rect 23406 11940 23430 11942
rect 23486 11940 23510 11942
rect 23566 11940 23572 11942
rect 23264 11931 23572 11940
rect 23676 11218 23704 12174
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23768 11694 23796 11834
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23264 10908 23572 10917
rect 23264 10906 23270 10908
rect 23326 10906 23350 10908
rect 23406 10906 23430 10908
rect 23486 10906 23510 10908
rect 23566 10906 23572 10908
rect 23326 10854 23328 10906
rect 23508 10854 23510 10906
rect 23264 10852 23270 10854
rect 23326 10852 23350 10854
rect 23406 10852 23430 10854
rect 23486 10852 23510 10854
rect 23566 10852 23572 10854
rect 23264 10843 23572 10852
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 22796 10220 22968 10248
rect 23020 10260 23072 10266
rect 22744 10202 22796 10208
rect 23020 10202 23072 10208
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22204 9846 22324 9874
rect 22008 8356 22060 8362
rect 22112 8350 22232 8378
rect 22008 8298 22060 8304
rect 22204 8294 22232 8350
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22112 7886 22140 8230
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 5234 22140 7686
rect 22204 7478 22232 7958
rect 22296 7478 22324 9846
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22388 6866 22416 10134
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22020 3194 22048 4082
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22112 3126 22140 4422
rect 22296 4282 22324 4966
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22296 3534 22324 3878
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21744 2746 21956 2774
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21744 2446 21772 2746
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 19524 2440 19576 2446
rect 16856 2382 16908 2388
rect 19430 2408 19486 2417
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 14936 1170 14964 2246
rect 14844 1142 14964 1170
rect 14844 800 14872 1142
rect 15488 800 15516 2246
rect 16132 870 16252 898
rect 16132 800 16160 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16224 762 16252 870
rect 16500 762 16528 2246
rect 16868 1306 16896 2382
rect 19340 2372 19392 2378
rect 19524 2382 19576 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 19430 2343 19486 2352
rect 19340 2314 19392 2320
rect 18052 2304 18104 2310
rect 18788 2304 18840 2310
rect 18052 2246 18104 2252
rect 18708 2264 18788 2292
rect 17077 2204 17385 2213
rect 17077 2202 17083 2204
rect 17139 2202 17163 2204
rect 17219 2202 17243 2204
rect 17299 2202 17323 2204
rect 17379 2202 17385 2204
rect 17139 2150 17141 2202
rect 17321 2150 17323 2202
rect 17077 2148 17083 2150
rect 17139 2148 17163 2150
rect 17219 2148 17243 2150
rect 17299 2148 17323 2150
rect 17379 2148 17385 2150
rect 17077 2139 17385 2148
rect 16776 1278 16896 1306
rect 16776 800 16804 1278
rect 18064 800 18092 2246
rect 18708 800 18736 2264
rect 18788 2246 18840 2252
rect 19352 1902 19380 2314
rect 19340 1896 19392 1902
rect 19340 1838 19392 1844
rect 19536 1306 19564 2382
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19996 1970 20024 2246
rect 19984 1964 20036 1970
rect 19984 1906 20036 1912
rect 20088 1306 20116 2382
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 19352 1278 19564 1306
rect 19996 1278 20116 1306
rect 19352 800 19380 1278
rect 19996 800 20024 1278
rect 21284 870 21404 898
rect 21284 800 21312 870
rect 16224 734 16528 762
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21376 762 21404 870
rect 21744 762 21772 2246
rect 21928 800 21956 2586
rect 22388 2038 22416 6054
rect 22376 2032 22428 2038
rect 22376 1974 22428 1980
rect 22480 1698 22508 9862
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22604 9276 22912 9285
rect 22604 9274 22610 9276
rect 22666 9274 22690 9276
rect 22746 9274 22770 9276
rect 22826 9274 22850 9276
rect 22906 9274 22912 9276
rect 22666 9222 22668 9274
rect 22848 9222 22850 9274
rect 22604 9220 22610 9222
rect 22666 9220 22690 9222
rect 22746 9220 22770 9222
rect 22826 9220 22850 9222
rect 22906 9220 22912 9222
rect 22604 9211 22912 9220
rect 22940 9178 22968 9454
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 22604 8188 22912 8197
rect 22604 8186 22610 8188
rect 22666 8186 22690 8188
rect 22746 8186 22770 8188
rect 22826 8186 22850 8188
rect 22906 8186 22912 8188
rect 22666 8134 22668 8186
rect 22848 8134 22850 8186
rect 22604 8132 22610 8134
rect 22666 8132 22690 8134
rect 22746 8132 22770 8134
rect 22826 8132 22850 8134
rect 22906 8132 22912 8134
rect 22604 8123 22912 8132
rect 22604 7100 22912 7109
rect 22604 7098 22610 7100
rect 22666 7098 22690 7100
rect 22746 7098 22770 7100
rect 22826 7098 22850 7100
rect 22906 7098 22912 7100
rect 22666 7046 22668 7098
rect 22848 7046 22850 7098
rect 22604 7044 22610 7046
rect 22666 7044 22690 7046
rect 22746 7044 22770 7046
rect 22826 7044 22850 7046
rect 22906 7044 22912 7046
rect 22604 7035 22912 7044
rect 22836 6112 22888 6118
rect 23032 6100 23060 9930
rect 23124 9722 23152 10610
rect 23676 10606 23704 11154
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23216 10266 23244 10406
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23676 10130 23704 10542
rect 23768 10198 23796 11630
rect 24044 11286 24072 12310
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24044 10470 24072 11222
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24044 10198 24072 10406
rect 23756 10192 23808 10198
rect 23756 10134 23808 10140
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23264 9820 23572 9829
rect 23264 9818 23270 9820
rect 23326 9818 23350 9820
rect 23406 9818 23430 9820
rect 23486 9818 23510 9820
rect 23566 9818 23572 9820
rect 23326 9766 23328 9818
rect 23508 9766 23510 9818
rect 23264 9764 23270 9766
rect 23326 9764 23350 9766
rect 23406 9764 23430 9766
rect 23486 9764 23510 9766
rect 23566 9764 23572 9766
rect 23264 9755 23572 9764
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23676 9654 23704 9862
rect 23768 9722 23796 10134
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23264 8732 23572 8741
rect 23264 8730 23270 8732
rect 23326 8730 23350 8732
rect 23406 8730 23430 8732
rect 23486 8730 23510 8732
rect 23566 8730 23572 8732
rect 23326 8678 23328 8730
rect 23508 8678 23510 8730
rect 23264 8676 23270 8678
rect 23326 8676 23350 8678
rect 23406 8676 23430 8678
rect 23486 8676 23510 8678
rect 23566 8676 23572 8678
rect 23264 8667 23572 8676
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23124 7478 23152 8230
rect 23264 7644 23572 7653
rect 23264 7642 23270 7644
rect 23326 7642 23350 7644
rect 23406 7642 23430 7644
rect 23486 7642 23510 7644
rect 23566 7642 23572 7644
rect 23326 7590 23328 7642
rect 23508 7590 23510 7642
rect 23264 7588 23270 7590
rect 23326 7588 23350 7590
rect 23406 7588 23430 7590
rect 23486 7588 23510 7590
rect 23566 7588 23572 7590
rect 23264 7579 23572 7588
rect 23112 7472 23164 7478
rect 23112 7414 23164 7420
rect 23264 6556 23572 6565
rect 23264 6554 23270 6556
rect 23326 6554 23350 6556
rect 23406 6554 23430 6556
rect 23486 6554 23510 6556
rect 23566 6554 23572 6556
rect 23326 6502 23328 6554
rect 23508 6502 23510 6554
rect 23264 6500 23270 6502
rect 23326 6500 23350 6502
rect 23406 6500 23430 6502
rect 23486 6500 23510 6502
rect 23566 6500 23572 6502
rect 23264 6491 23572 6500
rect 24136 6186 24164 17682
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24228 15162 24256 15302
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24320 10062 24348 23462
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24412 19446 24440 19654
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24504 18970 24532 25230
rect 24858 25191 24914 25200
rect 24964 21010 24992 25774
rect 25516 25498 25544 27911
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25792 25362 25820 28381
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25240 21622 25268 24142
rect 25412 24064 25464 24070
rect 25412 24006 25464 24012
rect 25424 23905 25452 24006
rect 25410 23896 25466 23905
rect 25410 23831 25466 23840
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24400 17808 24452 17814
rect 24400 17750 24452 17756
rect 24412 17338 24440 17750
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24412 12986 24440 15506
rect 24504 15502 24532 18022
rect 24688 17814 24716 19858
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24872 18970 24900 19790
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19514 25268 19654
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25410 19136 25466 19145
rect 25410 19071 25466 19080
rect 25424 18970 25452 19071
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25226 18864 25282 18873
rect 25226 18799 25282 18808
rect 25240 18766 25268 18799
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18358 24992 18566
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24872 17746 24900 18022
rect 25148 17882 25176 18702
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24504 14618 24532 14962
rect 24596 14890 24624 17002
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24688 15094 24716 16662
rect 24872 16590 24900 16934
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24964 15162 24992 16594
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 25056 16153 25084 16390
rect 25042 16144 25098 16153
rect 25042 16079 25098 16088
rect 25148 15994 25176 17478
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25240 16182 25268 16390
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25056 15966 25176 15994
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24596 14550 24624 14826
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24688 14346 24716 15030
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24688 14226 24716 14282
rect 24596 14198 24716 14226
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24504 13530 24532 13942
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24596 12918 24624 14198
rect 24780 13410 24808 14486
rect 24964 14414 24992 15098
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24872 13530 24900 14350
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24780 13382 24900 13410
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24688 12986 24716 13262
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24596 12306 24624 12854
rect 24872 12714 24900 13382
rect 25056 12714 25084 15966
rect 25240 15042 25268 15982
rect 25148 15014 25268 15042
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24872 12434 24900 12650
rect 24780 12406 24900 12434
rect 24780 12374 24808 12406
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 25148 11898 25176 15014
rect 25332 14906 25360 18022
rect 25516 15910 25544 23462
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25410 15736 25466 15745
rect 25410 15671 25412 15680
rect 25464 15671 25466 15680
rect 25412 15642 25464 15648
rect 25240 14878 25360 14906
rect 25240 14498 25268 14878
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25332 14618 25360 14758
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25240 14470 25360 14498
rect 25332 11898 25360 14470
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25424 13025 25452 13126
rect 25410 13016 25466 13025
rect 25410 12951 25466 12960
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11354 24440 11494
rect 24780 11354 24808 11698
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24412 10810 24440 10950
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24688 10674 24716 10950
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 24308 10056 24360 10062
rect 24964 10033 24992 10406
rect 25424 10305 25452 10406
rect 25410 10296 25466 10305
rect 25516 10266 25544 13806
rect 25608 13326 25636 23598
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25792 23225 25820 23462
rect 25778 23216 25834 23225
rect 25778 23151 25834 23160
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25688 17128 25740 17134
rect 25686 17096 25688 17105
rect 25740 17096 25742 17105
rect 25686 17031 25742 17040
rect 25686 13696 25742 13705
rect 25686 13631 25742 13640
rect 25700 13326 25728 13631
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25792 10674 25820 19314
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25410 10231 25466 10240
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 24308 9998 24360 10004
rect 24950 10024 25006 10033
rect 24950 9959 25006 9968
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9722 24900 9862
rect 24964 9722 24992 9959
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24504 9178 24532 9318
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24780 9042 24808 9454
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24124 6180 24176 6186
rect 24124 6122 24176 6128
rect 22888 6072 23060 6100
rect 22836 6054 22888 6060
rect 22604 6012 22912 6021
rect 22604 6010 22610 6012
rect 22666 6010 22690 6012
rect 22746 6010 22770 6012
rect 22826 6010 22850 6012
rect 22906 6010 22912 6012
rect 22666 5958 22668 6010
rect 22848 5958 22850 6010
rect 22604 5956 22610 5958
rect 22666 5956 22690 5958
rect 22746 5956 22770 5958
rect 22826 5956 22850 5958
rect 22906 5956 22912 5958
rect 22604 5947 22912 5956
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 22604 4924 22912 4933
rect 22604 4922 22610 4924
rect 22666 4922 22690 4924
rect 22746 4922 22770 4924
rect 22826 4922 22850 4924
rect 22906 4922 22912 4924
rect 22666 4870 22668 4922
rect 22848 4870 22850 4922
rect 22604 4868 22610 4870
rect 22666 4868 22690 4870
rect 22746 4868 22770 4870
rect 22826 4868 22850 4870
rect 22906 4868 22912 4870
rect 22604 4859 22912 4868
rect 22604 3836 22912 3845
rect 22604 3834 22610 3836
rect 22666 3834 22690 3836
rect 22746 3834 22770 3836
rect 22826 3834 22850 3836
rect 22906 3834 22912 3836
rect 22666 3782 22668 3834
rect 22848 3782 22850 3834
rect 22604 3780 22610 3782
rect 22666 3780 22690 3782
rect 22746 3780 22770 3782
rect 22826 3780 22850 3782
rect 22906 3780 22912 3782
rect 22604 3771 22912 3780
rect 23032 3534 23060 5170
rect 23124 4622 23152 5510
rect 23264 5468 23572 5477
rect 23264 5466 23270 5468
rect 23326 5466 23350 5468
rect 23406 5466 23430 5468
rect 23486 5466 23510 5468
rect 23566 5466 23572 5468
rect 23326 5414 23328 5466
rect 23508 5414 23510 5466
rect 23264 5412 23270 5414
rect 23326 5412 23350 5414
rect 23406 5412 23430 5414
rect 23486 5412 23510 5414
rect 23566 5412 23572 5414
rect 23264 5403 23572 5412
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3126 22876 3334
rect 23124 3126 23152 4558
rect 23264 4380 23572 4389
rect 23264 4378 23270 4380
rect 23326 4378 23350 4380
rect 23406 4378 23430 4380
rect 23486 4378 23510 4380
rect 23566 4378 23572 4380
rect 23326 4326 23328 4378
rect 23508 4326 23510 4378
rect 23264 4324 23270 4326
rect 23326 4324 23350 4326
rect 23406 4324 23430 4326
rect 23486 4324 23510 4326
rect 23566 4324 23572 4326
rect 23264 4315 23572 4324
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23676 3738 23704 3878
rect 24780 3738 24808 8774
rect 24872 3738 24900 9522
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 25240 8362 25268 8978
rect 25332 8566 25360 9318
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24964 3942 24992 7686
rect 25240 4622 25268 8298
rect 25516 6322 25544 10202
rect 25884 8362 25912 26318
rect 26436 25906 26464 28381
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26148 25220 26200 25226
rect 26148 25162 26200 25168
rect 25964 22568 26016 22574
rect 25962 22536 25964 22545
rect 26016 22536 26018 22545
rect 25962 22471 26018 22480
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25976 21865 26004 21898
rect 25962 21856 26018 21865
rect 25962 21791 26018 21800
rect 25964 20732 26016 20738
rect 25964 20674 26016 20680
rect 25976 20505 26004 20674
rect 25962 20496 26018 20505
rect 25962 20431 26018 20440
rect 25964 19984 26016 19990
rect 25964 19926 26016 19932
rect 25976 19825 26004 19926
rect 26056 19848 26108 19854
rect 25962 19816 26018 19825
rect 26056 19790 26108 19796
rect 25962 19751 26018 19760
rect 25962 18456 26018 18465
rect 25962 18391 26018 18400
rect 25976 18358 26004 18391
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25964 17060 26016 17066
rect 25964 17002 26016 17008
rect 25976 16425 26004 17002
rect 25962 16416 26018 16425
rect 25962 16351 26018 16360
rect 25964 14544 26016 14550
rect 25964 14486 26016 14492
rect 25976 14385 26004 14486
rect 25962 14376 26018 14385
rect 25962 14311 26018 14320
rect 26068 14226 26096 19790
rect 26160 16250 26188 25162
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26252 15502 26280 22374
rect 26332 21072 26384 21078
rect 26332 21014 26384 21020
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 25976 14198 26096 14226
rect 25976 12170 26004 14198
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 26068 12345 26096 12786
rect 26344 12753 26372 21014
rect 26330 12744 26386 12753
rect 26330 12679 26386 12688
rect 26054 12336 26110 12345
rect 26054 12271 26110 12280
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25976 10985 26004 11018
rect 25962 10976 26018 10985
rect 25962 10911 26018 10920
rect 25964 9784 26016 9790
rect 25964 9726 26016 9732
rect 25976 9625 26004 9726
rect 25962 9616 26018 9625
rect 25962 9551 26018 9560
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25962 8256 26018 8265
rect 25962 8191 26018 8200
rect 25976 7886 26004 8191
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25700 7585 25728 7686
rect 25686 7576 25742 7585
rect 25686 7511 25742 7520
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 25976 6905 26004 6938
rect 25962 6896 26018 6905
rect 25962 6831 26018 6840
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25410 6216 25466 6225
rect 25410 6151 25412 6160
rect 25464 6151 25466 6160
rect 25412 6122 25464 6128
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4865 25452 4966
rect 25410 4856 25466 4865
rect 25410 4791 25466 4800
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25424 4185 25452 4422
rect 25410 4176 25466 4185
rect 25410 4111 25466 4120
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 23264 3292 23572 3301
rect 23264 3290 23270 3292
rect 23326 3290 23350 3292
rect 23406 3290 23430 3292
rect 23486 3290 23510 3292
rect 23566 3290 23572 3292
rect 23326 3238 23328 3290
rect 23508 3238 23510 3290
rect 23264 3236 23270 3238
rect 23326 3236 23350 3238
rect 23406 3236 23430 3238
rect 23486 3236 23510 3238
rect 23566 3236 23572 3238
rect 23264 3227 23572 3236
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 24688 3058 24716 3470
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24676 3052 24728 3058
rect 24676 2994 24728 3000
rect 22604 2748 22912 2757
rect 22604 2746 22610 2748
rect 22666 2746 22690 2748
rect 22746 2746 22770 2748
rect 22826 2746 22850 2748
rect 22906 2746 22912 2748
rect 22666 2694 22668 2746
rect 22848 2694 22850 2746
rect 22604 2692 22610 2694
rect 22666 2692 22690 2694
rect 22746 2692 22770 2694
rect 22826 2692 22850 2694
rect 22906 2692 22912 2694
rect 22604 2683 22912 2692
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 22468 1692 22520 1698
rect 22468 1634 22520 1640
rect 22664 1170 22692 2382
rect 22940 2106 22968 2382
rect 23264 2204 23572 2213
rect 23264 2202 23270 2204
rect 23326 2202 23350 2204
rect 23406 2202 23430 2204
rect 23486 2202 23510 2204
rect 23566 2202 23572 2204
rect 23326 2150 23328 2202
rect 23508 2150 23510 2202
rect 23264 2148 23270 2150
rect 23326 2148 23350 2150
rect 23406 2148 23430 2150
rect 23486 2148 23510 2150
rect 23566 2148 23572 2150
rect 23264 2139 23572 2148
rect 22928 2100 22980 2106
rect 22928 2042 22980 2048
rect 23952 1306 23980 2382
rect 24596 1562 24624 2994
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 24584 1556 24636 1562
rect 24584 1498 24636 1504
rect 24688 1465 24716 2858
rect 24872 2446 24900 3538
rect 24952 3528 25004 3534
rect 25964 3528 26016 3534
rect 24952 3470 25004 3476
rect 25962 3496 25964 3505
rect 26016 3496 26018 3505
rect 24964 2774 24992 3470
rect 25872 3460 25924 3466
rect 25962 3431 26018 3440
rect 25872 3402 25924 3408
rect 25136 2848 25188 2854
rect 25134 2816 25136 2825
rect 25188 2816 25190 2825
rect 24964 2746 25084 2774
rect 25134 2751 25190 2760
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24860 2304 24912 2310
rect 24780 2264 24860 2292
rect 24674 1456 24730 1465
rect 24674 1391 24730 1400
rect 22572 1142 22692 1170
rect 23860 1278 23980 1306
rect 22572 800 22600 1142
rect 23860 800 23888 1278
rect 24504 870 24624 898
rect 24504 800 24532 870
rect 21376 734 21772 762
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 24596 762 24624 870
rect 24780 762 24808 2264
rect 24860 2246 24912 2252
rect 25056 921 25084 2746
rect 25228 2304 25280 2310
rect 25148 2264 25228 2292
rect 25042 912 25098 921
rect 25042 847 25098 856
rect 25148 800 25176 2264
rect 25228 2246 25280 2252
rect 25780 1556 25832 1562
rect 25780 1498 25832 1504
rect 25792 800 25820 1498
rect 24596 734 24808 762
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 25884 105 25912 3402
rect 25870 96 25926 105
rect 25870 31 25926 40
<< via2 >>
rect 1582 28600 1638 28656
rect 1398 26968 1454 27024
rect 1030 25880 1086 25936
rect 2870 26560 2926 26616
rect 1030 25236 1032 25256
rect 1032 25236 1084 25256
rect 1084 25236 1086 25256
rect 1030 25200 1086 25236
rect 938 23840 994 23896
rect 1582 23588 1638 23624
rect 1582 23568 1584 23588
rect 1584 23568 1636 23588
rect 1636 23568 1638 23588
rect 1398 23432 1454 23488
rect 938 22480 994 22536
rect 938 21120 994 21176
rect 1398 20576 1454 20632
rect 1582 19508 1638 19544
rect 1582 19488 1584 19508
rect 1584 19488 1636 19508
rect 1636 19488 1638 19508
rect 1490 19372 1546 19408
rect 1490 19352 1492 19372
rect 1492 19352 1544 19372
rect 1544 19352 1546 19372
rect 1490 18284 1546 18320
rect 1490 18264 1492 18284
rect 1492 18264 1544 18284
rect 1544 18264 1546 18284
rect 938 17076 940 17096
rect 940 17076 992 17096
rect 992 17076 994 17096
rect 938 17040 994 17076
rect 1398 16496 1454 16552
rect 938 15680 994 15736
rect 938 14356 940 14376
rect 940 14356 992 14376
rect 992 14356 994 14376
rect 938 14320 994 14356
rect 1398 13640 1454 13696
rect 938 12960 994 13016
rect 1582 17856 1638 17912
rect 1582 17060 1638 17096
rect 1582 17040 1584 17060
rect 1584 17040 1636 17060
rect 1636 17040 1638 17060
rect 2410 21392 2466 21448
rect 1950 19216 2006 19272
rect 1858 16088 1914 16144
rect 1766 15408 1822 15464
rect 938 11600 994 11656
rect 938 10240 994 10296
rect 1582 10956 1584 10976
rect 1584 10956 1636 10976
rect 1636 10956 1638 10976
rect 1582 10920 1638 10956
rect 1490 10668 1546 10704
rect 1490 10648 1492 10668
rect 1492 10648 1544 10668
rect 1544 10648 1546 10668
rect 1674 10104 1730 10160
rect 938 9560 994 9616
rect 1674 8200 1730 8256
rect 938 7540 994 7576
rect 938 7520 940 7540
rect 940 7520 992 7540
rect 992 7520 994 7540
rect 2686 20440 2742 20496
rect 2962 20340 2964 20360
rect 2964 20340 3016 20360
rect 3016 20340 3018 20360
rect 2962 20304 3018 20340
rect 2134 9968 2190 10024
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 938 4800 994 4856
rect 1582 4528 1638 4584
rect 938 4120 994 4176
rect 1030 3476 1032 3496
rect 1032 3476 1084 3496
rect 1084 3476 1086 3496
rect 1030 3440 1086 3476
rect 4049 26682 4105 26684
rect 4129 26682 4185 26684
rect 4209 26682 4265 26684
rect 4289 26682 4345 26684
rect 4049 26630 4095 26682
rect 4095 26630 4105 26682
rect 4129 26630 4159 26682
rect 4159 26630 4171 26682
rect 4171 26630 4185 26682
rect 4209 26630 4223 26682
rect 4223 26630 4235 26682
rect 4235 26630 4265 26682
rect 4289 26630 4299 26682
rect 4299 26630 4345 26682
rect 4049 26628 4105 26630
rect 4129 26628 4185 26630
rect 4209 26628 4265 26630
rect 4289 26628 4345 26630
rect 4709 26138 4765 26140
rect 4789 26138 4845 26140
rect 4869 26138 4925 26140
rect 4949 26138 5005 26140
rect 4709 26086 4755 26138
rect 4755 26086 4765 26138
rect 4789 26086 4819 26138
rect 4819 26086 4831 26138
rect 4831 26086 4845 26138
rect 4869 26086 4883 26138
rect 4883 26086 4895 26138
rect 4895 26086 4925 26138
rect 4949 26086 4959 26138
rect 4959 26086 5005 26138
rect 4709 26084 4765 26086
rect 4789 26084 4845 26086
rect 4869 26084 4925 26086
rect 4949 26084 5005 26086
rect 4049 25594 4105 25596
rect 4129 25594 4185 25596
rect 4209 25594 4265 25596
rect 4289 25594 4345 25596
rect 4049 25542 4095 25594
rect 4095 25542 4105 25594
rect 4129 25542 4159 25594
rect 4159 25542 4171 25594
rect 4171 25542 4185 25594
rect 4209 25542 4223 25594
rect 4223 25542 4235 25594
rect 4235 25542 4265 25594
rect 4289 25542 4299 25594
rect 4299 25542 4345 25594
rect 4049 25540 4105 25542
rect 4129 25540 4185 25542
rect 4209 25540 4265 25542
rect 4289 25540 4345 25542
rect 4709 25050 4765 25052
rect 4789 25050 4845 25052
rect 4869 25050 4925 25052
rect 4949 25050 5005 25052
rect 4709 24998 4755 25050
rect 4755 24998 4765 25050
rect 4789 24998 4819 25050
rect 4819 24998 4831 25050
rect 4831 24998 4845 25050
rect 4869 24998 4883 25050
rect 4883 24998 4895 25050
rect 4895 24998 4925 25050
rect 4949 24998 4959 25050
rect 4959 24998 5005 25050
rect 4709 24996 4765 24998
rect 4789 24996 4845 24998
rect 4869 24996 4925 24998
rect 4949 24996 5005 24998
rect 4049 24506 4105 24508
rect 4129 24506 4185 24508
rect 4209 24506 4265 24508
rect 4289 24506 4345 24508
rect 4049 24454 4095 24506
rect 4095 24454 4105 24506
rect 4129 24454 4159 24506
rect 4159 24454 4171 24506
rect 4171 24454 4185 24506
rect 4209 24454 4223 24506
rect 4223 24454 4235 24506
rect 4235 24454 4265 24506
rect 4289 24454 4299 24506
rect 4299 24454 4345 24506
rect 4049 24452 4105 24454
rect 4129 24452 4185 24454
rect 4209 24452 4265 24454
rect 4289 24452 4345 24454
rect 4709 23962 4765 23964
rect 4789 23962 4845 23964
rect 4869 23962 4925 23964
rect 4949 23962 5005 23964
rect 4709 23910 4755 23962
rect 4755 23910 4765 23962
rect 4789 23910 4819 23962
rect 4819 23910 4831 23962
rect 4831 23910 4845 23962
rect 4869 23910 4883 23962
rect 4883 23910 4895 23962
rect 4895 23910 4925 23962
rect 4949 23910 4959 23962
rect 4959 23910 5005 23962
rect 4709 23908 4765 23910
rect 4789 23908 4845 23910
rect 4869 23908 4925 23910
rect 4949 23908 5005 23910
rect 4049 23418 4105 23420
rect 4129 23418 4185 23420
rect 4209 23418 4265 23420
rect 4289 23418 4345 23420
rect 4049 23366 4095 23418
rect 4095 23366 4105 23418
rect 4129 23366 4159 23418
rect 4159 23366 4171 23418
rect 4171 23366 4185 23418
rect 4209 23366 4223 23418
rect 4223 23366 4235 23418
rect 4235 23366 4265 23418
rect 4289 23366 4299 23418
rect 4299 23366 4345 23418
rect 4049 23364 4105 23366
rect 4129 23364 4185 23366
rect 4209 23364 4265 23366
rect 4289 23364 4345 23366
rect 4049 22330 4105 22332
rect 4129 22330 4185 22332
rect 4209 22330 4265 22332
rect 4289 22330 4345 22332
rect 4049 22278 4095 22330
rect 4095 22278 4105 22330
rect 4129 22278 4159 22330
rect 4159 22278 4171 22330
rect 4171 22278 4185 22330
rect 4209 22278 4223 22330
rect 4223 22278 4235 22330
rect 4235 22278 4265 22330
rect 4289 22278 4299 22330
rect 4299 22278 4345 22330
rect 4049 22276 4105 22278
rect 4129 22276 4185 22278
rect 4209 22276 4265 22278
rect 4289 22276 4345 22278
rect 4049 21242 4105 21244
rect 4129 21242 4185 21244
rect 4209 21242 4265 21244
rect 4289 21242 4345 21244
rect 4049 21190 4095 21242
rect 4095 21190 4105 21242
rect 4129 21190 4159 21242
rect 4159 21190 4171 21242
rect 4171 21190 4185 21242
rect 4209 21190 4223 21242
rect 4223 21190 4235 21242
rect 4235 21190 4265 21242
rect 4289 21190 4299 21242
rect 4299 21190 4345 21242
rect 4049 21188 4105 21190
rect 4129 21188 4185 21190
rect 4209 21188 4265 21190
rect 4289 21188 4345 21190
rect 4709 22874 4765 22876
rect 4789 22874 4845 22876
rect 4869 22874 4925 22876
rect 4949 22874 5005 22876
rect 4709 22822 4755 22874
rect 4755 22822 4765 22874
rect 4789 22822 4819 22874
rect 4819 22822 4831 22874
rect 4831 22822 4845 22874
rect 4869 22822 4883 22874
rect 4883 22822 4895 22874
rect 4895 22822 4925 22874
rect 4949 22822 4959 22874
rect 4959 22822 5005 22874
rect 4709 22820 4765 22822
rect 4789 22820 4845 22822
rect 4869 22820 4925 22822
rect 4949 22820 5005 22822
rect 4709 21786 4765 21788
rect 4789 21786 4845 21788
rect 4869 21786 4925 21788
rect 4949 21786 5005 21788
rect 4709 21734 4755 21786
rect 4755 21734 4765 21786
rect 4789 21734 4819 21786
rect 4819 21734 4831 21786
rect 4831 21734 4845 21786
rect 4869 21734 4883 21786
rect 4883 21734 4895 21786
rect 4895 21734 4925 21786
rect 4949 21734 4959 21786
rect 4959 21734 5005 21786
rect 4709 21732 4765 21734
rect 4789 21732 4845 21734
rect 4869 21732 4925 21734
rect 4949 21732 5005 21734
rect 4049 20154 4105 20156
rect 4129 20154 4185 20156
rect 4209 20154 4265 20156
rect 4289 20154 4345 20156
rect 4049 20102 4095 20154
rect 4095 20102 4105 20154
rect 4129 20102 4159 20154
rect 4159 20102 4171 20154
rect 4171 20102 4185 20154
rect 4209 20102 4223 20154
rect 4223 20102 4235 20154
rect 4235 20102 4265 20154
rect 4289 20102 4299 20154
rect 4299 20102 4345 20154
rect 4049 20100 4105 20102
rect 4129 20100 4185 20102
rect 4209 20100 4265 20102
rect 4289 20100 4345 20102
rect 4250 19916 4306 19952
rect 4250 19896 4252 19916
rect 4252 19896 4304 19916
rect 4304 19896 4306 19916
rect 4709 20698 4765 20700
rect 4789 20698 4845 20700
rect 4869 20698 4925 20700
rect 4949 20698 5005 20700
rect 4709 20646 4755 20698
rect 4755 20646 4765 20698
rect 4789 20646 4819 20698
rect 4819 20646 4831 20698
rect 4831 20646 4845 20698
rect 4869 20646 4883 20698
rect 4883 20646 4895 20698
rect 4895 20646 4925 20698
rect 4949 20646 4959 20698
rect 4959 20646 5005 20698
rect 4709 20644 4765 20646
rect 4789 20644 4845 20646
rect 4869 20644 4925 20646
rect 4949 20644 5005 20646
rect 4049 19066 4105 19068
rect 4129 19066 4185 19068
rect 4209 19066 4265 19068
rect 4289 19066 4345 19068
rect 4049 19014 4095 19066
rect 4095 19014 4105 19066
rect 4129 19014 4159 19066
rect 4159 19014 4171 19066
rect 4171 19014 4185 19066
rect 4209 19014 4223 19066
rect 4223 19014 4235 19066
rect 4235 19014 4265 19066
rect 4289 19014 4299 19066
rect 4299 19014 4345 19066
rect 4049 19012 4105 19014
rect 4129 19012 4185 19014
rect 4209 19012 4265 19014
rect 4289 19012 4345 19014
rect 4158 18808 4214 18864
rect 4250 18672 4306 18728
rect 4526 19252 4528 19272
rect 4528 19252 4580 19272
rect 4580 19252 4582 19272
rect 4526 19216 4582 19252
rect 4709 19610 4765 19612
rect 4789 19610 4845 19612
rect 4869 19610 4925 19612
rect 4949 19610 5005 19612
rect 4709 19558 4755 19610
rect 4755 19558 4765 19610
rect 4789 19558 4819 19610
rect 4819 19558 4831 19610
rect 4831 19558 4845 19610
rect 4869 19558 4883 19610
rect 4883 19558 4895 19610
rect 4895 19558 4925 19610
rect 4949 19558 4959 19610
rect 4959 19558 5005 19610
rect 4709 19556 4765 19558
rect 4789 19556 4845 19558
rect 4869 19556 4925 19558
rect 4949 19556 5005 19558
rect 10236 26682 10292 26684
rect 10316 26682 10372 26684
rect 10396 26682 10452 26684
rect 10476 26682 10532 26684
rect 10236 26630 10282 26682
rect 10282 26630 10292 26682
rect 10316 26630 10346 26682
rect 10346 26630 10358 26682
rect 10358 26630 10372 26682
rect 10396 26630 10410 26682
rect 10410 26630 10422 26682
rect 10422 26630 10452 26682
rect 10476 26630 10486 26682
rect 10486 26630 10532 26682
rect 10236 26628 10292 26630
rect 10316 26628 10372 26630
rect 10396 26628 10452 26630
rect 10476 26628 10532 26630
rect 4802 18944 4858 19000
rect 4802 18808 4858 18864
rect 4049 17978 4105 17980
rect 4129 17978 4185 17980
rect 4209 17978 4265 17980
rect 4289 17978 4345 17980
rect 4049 17926 4095 17978
rect 4095 17926 4105 17978
rect 4129 17926 4159 17978
rect 4159 17926 4171 17978
rect 4171 17926 4185 17978
rect 4209 17926 4223 17978
rect 4223 17926 4235 17978
rect 4235 17926 4265 17978
rect 4289 17926 4299 17978
rect 4299 17926 4345 17978
rect 4049 17924 4105 17926
rect 4129 17924 4185 17926
rect 4209 17924 4265 17926
rect 4289 17924 4345 17926
rect 4709 18522 4765 18524
rect 4789 18522 4845 18524
rect 4869 18522 4925 18524
rect 4949 18522 5005 18524
rect 4709 18470 4755 18522
rect 4755 18470 4765 18522
rect 4789 18470 4819 18522
rect 4819 18470 4831 18522
rect 4831 18470 4845 18522
rect 4869 18470 4883 18522
rect 4883 18470 4895 18522
rect 4895 18470 4925 18522
rect 4949 18470 4959 18522
rect 4959 18470 5005 18522
rect 4709 18468 4765 18470
rect 4789 18468 4845 18470
rect 4869 18468 4925 18470
rect 4949 18468 5005 18470
rect 4709 17434 4765 17436
rect 4789 17434 4845 17436
rect 4869 17434 4925 17436
rect 4949 17434 5005 17436
rect 4709 17382 4755 17434
rect 4755 17382 4765 17434
rect 4789 17382 4819 17434
rect 4819 17382 4831 17434
rect 4831 17382 4845 17434
rect 4869 17382 4883 17434
rect 4883 17382 4895 17434
rect 4895 17382 4925 17434
rect 4949 17382 4959 17434
rect 4959 17382 5005 17434
rect 4709 17380 4765 17382
rect 4789 17380 4845 17382
rect 4869 17380 4925 17382
rect 4949 17380 5005 17382
rect 4049 16890 4105 16892
rect 4129 16890 4185 16892
rect 4209 16890 4265 16892
rect 4289 16890 4345 16892
rect 4049 16838 4095 16890
rect 4095 16838 4105 16890
rect 4129 16838 4159 16890
rect 4159 16838 4171 16890
rect 4171 16838 4185 16890
rect 4209 16838 4223 16890
rect 4223 16838 4235 16890
rect 4235 16838 4265 16890
rect 4289 16838 4299 16890
rect 4299 16838 4345 16890
rect 4049 16836 4105 16838
rect 4129 16836 4185 16838
rect 4209 16836 4265 16838
rect 4289 16836 4345 16838
rect 4709 16346 4765 16348
rect 4789 16346 4845 16348
rect 4869 16346 4925 16348
rect 4949 16346 5005 16348
rect 4709 16294 4755 16346
rect 4755 16294 4765 16346
rect 4789 16294 4819 16346
rect 4819 16294 4831 16346
rect 4831 16294 4845 16346
rect 4869 16294 4883 16346
rect 4883 16294 4895 16346
rect 4895 16294 4925 16346
rect 4949 16294 4959 16346
rect 4959 16294 5005 16346
rect 4709 16292 4765 16294
rect 4789 16292 4845 16294
rect 4869 16292 4925 16294
rect 4949 16292 5005 16294
rect 4049 15802 4105 15804
rect 4129 15802 4185 15804
rect 4209 15802 4265 15804
rect 4289 15802 4345 15804
rect 4049 15750 4095 15802
rect 4095 15750 4105 15802
rect 4129 15750 4159 15802
rect 4159 15750 4171 15802
rect 4171 15750 4185 15802
rect 4209 15750 4223 15802
rect 4223 15750 4235 15802
rect 4235 15750 4265 15802
rect 4289 15750 4299 15802
rect 4299 15750 4345 15802
rect 4049 15748 4105 15750
rect 4129 15748 4185 15750
rect 4209 15748 4265 15750
rect 4289 15748 4345 15750
rect 4709 15258 4765 15260
rect 4789 15258 4845 15260
rect 4869 15258 4925 15260
rect 4949 15258 5005 15260
rect 4709 15206 4755 15258
rect 4755 15206 4765 15258
rect 4789 15206 4819 15258
rect 4819 15206 4831 15258
rect 4831 15206 4845 15258
rect 4869 15206 4883 15258
rect 4883 15206 4895 15258
rect 4895 15206 4925 15258
rect 4949 15206 4959 15258
rect 4959 15206 5005 15258
rect 4709 15204 4765 15206
rect 4789 15204 4845 15206
rect 4869 15204 4925 15206
rect 4949 15204 5005 15206
rect 4049 14714 4105 14716
rect 4129 14714 4185 14716
rect 4209 14714 4265 14716
rect 4289 14714 4345 14716
rect 4049 14662 4095 14714
rect 4095 14662 4105 14714
rect 4129 14662 4159 14714
rect 4159 14662 4171 14714
rect 4171 14662 4185 14714
rect 4209 14662 4223 14714
rect 4223 14662 4235 14714
rect 4235 14662 4265 14714
rect 4289 14662 4299 14714
rect 4299 14662 4345 14714
rect 4049 14660 4105 14662
rect 4129 14660 4185 14662
rect 4209 14660 4265 14662
rect 4289 14660 4345 14662
rect 4049 13626 4105 13628
rect 4129 13626 4185 13628
rect 4209 13626 4265 13628
rect 4289 13626 4345 13628
rect 4049 13574 4095 13626
rect 4095 13574 4105 13626
rect 4129 13574 4159 13626
rect 4159 13574 4171 13626
rect 4171 13574 4185 13626
rect 4209 13574 4223 13626
rect 4223 13574 4235 13626
rect 4235 13574 4265 13626
rect 4289 13574 4299 13626
rect 4299 13574 4345 13626
rect 4049 13572 4105 13574
rect 4129 13572 4185 13574
rect 4209 13572 4265 13574
rect 4289 13572 4345 13574
rect 4342 13232 4398 13288
rect 4709 14170 4765 14172
rect 4789 14170 4845 14172
rect 4869 14170 4925 14172
rect 4949 14170 5005 14172
rect 4709 14118 4755 14170
rect 4755 14118 4765 14170
rect 4789 14118 4819 14170
rect 4819 14118 4831 14170
rect 4831 14118 4845 14170
rect 4869 14118 4883 14170
rect 4883 14118 4895 14170
rect 4895 14118 4925 14170
rect 4949 14118 4959 14170
rect 4959 14118 5005 14170
rect 4709 14116 4765 14118
rect 4789 14116 4845 14118
rect 4869 14116 4925 14118
rect 4949 14116 5005 14118
rect 5262 18844 5264 18864
rect 5264 18844 5316 18864
rect 5316 18844 5318 18864
rect 5262 18808 5318 18844
rect 5262 17856 5318 17912
rect 5446 17720 5502 17776
rect 5538 17584 5594 17640
rect 4049 12538 4105 12540
rect 4129 12538 4185 12540
rect 4209 12538 4265 12540
rect 4289 12538 4345 12540
rect 4049 12486 4095 12538
rect 4095 12486 4105 12538
rect 4129 12486 4159 12538
rect 4159 12486 4171 12538
rect 4171 12486 4185 12538
rect 4209 12486 4223 12538
rect 4223 12486 4235 12538
rect 4235 12486 4265 12538
rect 4289 12486 4299 12538
rect 4299 12486 4345 12538
rect 4049 12484 4105 12486
rect 4129 12484 4185 12486
rect 4209 12484 4265 12486
rect 4289 12484 4345 12486
rect 4709 13082 4765 13084
rect 4789 13082 4845 13084
rect 4869 13082 4925 13084
rect 4949 13082 5005 13084
rect 4709 13030 4755 13082
rect 4755 13030 4765 13082
rect 4789 13030 4819 13082
rect 4819 13030 4831 13082
rect 4831 13030 4845 13082
rect 4869 13030 4883 13082
rect 4883 13030 4895 13082
rect 4895 13030 4925 13082
rect 4949 13030 4959 13082
rect 4959 13030 5005 13082
rect 4709 13028 4765 13030
rect 4789 13028 4845 13030
rect 4869 13028 4925 13030
rect 4949 13028 5005 13030
rect 4049 11450 4105 11452
rect 4129 11450 4185 11452
rect 4209 11450 4265 11452
rect 4289 11450 4345 11452
rect 4049 11398 4095 11450
rect 4095 11398 4105 11450
rect 4129 11398 4159 11450
rect 4159 11398 4171 11450
rect 4171 11398 4185 11450
rect 4209 11398 4223 11450
rect 4223 11398 4235 11450
rect 4235 11398 4265 11450
rect 4289 11398 4299 11450
rect 4299 11398 4345 11450
rect 4049 11396 4105 11398
rect 4129 11396 4185 11398
rect 4209 11396 4265 11398
rect 4289 11396 4345 11398
rect 4049 10362 4105 10364
rect 4129 10362 4185 10364
rect 4209 10362 4265 10364
rect 4289 10362 4345 10364
rect 4049 10310 4095 10362
rect 4095 10310 4105 10362
rect 4129 10310 4159 10362
rect 4159 10310 4171 10362
rect 4171 10310 4185 10362
rect 4209 10310 4223 10362
rect 4223 10310 4235 10362
rect 4235 10310 4265 10362
rect 4289 10310 4299 10362
rect 4299 10310 4345 10362
rect 4049 10308 4105 10310
rect 4129 10308 4185 10310
rect 4209 10308 4265 10310
rect 4289 10308 4345 10310
rect 5446 16516 5502 16552
rect 5446 16496 5448 16516
rect 5448 16496 5500 16516
rect 5500 16496 5502 16516
rect 4709 11994 4765 11996
rect 4789 11994 4845 11996
rect 4869 11994 4925 11996
rect 4949 11994 5005 11996
rect 4709 11942 4755 11994
rect 4755 11942 4765 11994
rect 4789 11942 4819 11994
rect 4819 11942 4831 11994
rect 4831 11942 4845 11994
rect 4869 11942 4883 11994
rect 4883 11942 4895 11994
rect 4895 11942 4925 11994
rect 4949 11942 4959 11994
rect 4959 11942 5005 11994
rect 4709 11940 4765 11942
rect 4789 11940 4845 11942
rect 4869 11940 4925 11942
rect 4949 11940 5005 11942
rect 4709 10906 4765 10908
rect 4789 10906 4845 10908
rect 4869 10906 4925 10908
rect 4949 10906 5005 10908
rect 4709 10854 4755 10906
rect 4755 10854 4765 10906
rect 4789 10854 4819 10906
rect 4819 10854 4831 10906
rect 4831 10854 4845 10906
rect 4869 10854 4883 10906
rect 4883 10854 4895 10906
rect 4895 10854 4925 10906
rect 4949 10854 4959 10906
rect 4959 10854 5005 10906
rect 4709 10852 4765 10854
rect 4789 10852 4845 10854
rect 4869 10852 4925 10854
rect 4949 10852 5005 10854
rect 5078 10512 5134 10568
rect 4709 9818 4765 9820
rect 4789 9818 4845 9820
rect 4869 9818 4925 9820
rect 4949 9818 5005 9820
rect 4709 9766 4755 9818
rect 4755 9766 4765 9818
rect 4789 9766 4819 9818
rect 4819 9766 4831 9818
rect 4831 9766 4845 9818
rect 4869 9766 4883 9818
rect 4883 9766 4895 9818
rect 4895 9766 4925 9818
rect 4949 9766 4959 9818
rect 4959 9766 5005 9818
rect 4709 9764 4765 9766
rect 4789 9764 4845 9766
rect 4869 9764 4925 9766
rect 4949 9764 5005 9766
rect 4250 9580 4306 9616
rect 4250 9560 4252 9580
rect 4252 9560 4304 9580
rect 4304 9560 4306 9580
rect 4049 9274 4105 9276
rect 4129 9274 4185 9276
rect 4209 9274 4265 9276
rect 4289 9274 4345 9276
rect 4049 9222 4095 9274
rect 4095 9222 4105 9274
rect 4129 9222 4159 9274
rect 4159 9222 4171 9274
rect 4171 9222 4185 9274
rect 4209 9222 4223 9274
rect 4223 9222 4235 9274
rect 4235 9222 4265 9274
rect 4289 9222 4299 9274
rect 4299 9222 4345 9274
rect 4049 9220 4105 9222
rect 4129 9220 4185 9222
rect 4209 9220 4265 9222
rect 4289 9220 4345 9222
rect 4709 8730 4765 8732
rect 4789 8730 4845 8732
rect 4869 8730 4925 8732
rect 4949 8730 5005 8732
rect 4709 8678 4755 8730
rect 4755 8678 4765 8730
rect 4789 8678 4819 8730
rect 4819 8678 4831 8730
rect 4831 8678 4845 8730
rect 4869 8678 4883 8730
rect 4883 8678 4895 8730
rect 4895 8678 4925 8730
rect 4949 8678 4959 8730
rect 4959 8678 5005 8730
rect 4709 8676 4765 8678
rect 4789 8676 4845 8678
rect 4869 8676 4925 8678
rect 4949 8676 5005 8678
rect 4049 8186 4105 8188
rect 4129 8186 4185 8188
rect 4209 8186 4265 8188
rect 4289 8186 4345 8188
rect 4049 8134 4095 8186
rect 4095 8134 4105 8186
rect 4129 8134 4159 8186
rect 4159 8134 4171 8186
rect 4171 8134 4185 8186
rect 4209 8134 4223 8186
rect 4223 8134 4235 8186
rect 4235 8134 4265 8186
rect 4289 8134 4299 8186
rect 4299 8134 4345 8186
rect 4049 8132 4105 8134
rect 4129 8132 4185 8134
rect 4209 8132 4265 8134
rect 4289 8132 4345 8134
rect 2778 6840 2834 6896
rect 4049 7098 4105 7100
rect 4129 7098 4185 7100
rect 4209 7098 4265 7100
rect 4289 7098 4345 7100
rect 4049 7046 4095 7098
rect 4095 7046 4105 7098
rect 4129 7046 4159 7098
rect 4159 7046 4171 7098
rect 4171 7046 4185 7098
rect 4209 7046 4223 7098
rect 4223 7046 4235 7098
rect 4235 7046 4265 7098
rect 4289 7046 4299 7098
rect 4299 7046 4345 7098
rect 4049 7044 4105 7046
rect 4129 7044 4185 7046
rect 4209 7044 4265 7046
rect 4289 7044 4345 7046
rect 4049 6010 4105 6012
rect 4129 6010 4185 6012
rect 4209 6010 4265 6012
rect 4289 6010 4345 6012
rect 4049 5958 4095 6010
rect 4095 5958 4105 6010
rect 4129 5958 4159 6010
rect 4159 5958 4171 6010
rect 4171 5958 4185 6010
rect 4209 5958 4223 6010
rect 4223 5958 4235 6010
rect 4235 5958 4265 6010
rect 4289 5958 4299 6010
rect 4299 5958 4345 6010
rect 4049 5956 4105 5958
rect 4129 5956 4185 5958
rect 4209 5956 4265 5958
rect 4289 5956 4345 5958
rect 4709 7642 4765 7644
rect 4789 7642 4845 7644
rect 4869 7642 4925 7644
rect 4949 7642 5005 7644
rect 4709 7590 4755 7642
rect 4755 7590 4765 7642
rect 4789 7590 4819 7642
rect 4819 7590 4831 7642
rect 4831 7590 4845 7642
rect 4869 7590 4883 7642
rect 4883 7590 4895 7642
rect 4895 7590 4925 7642
rect 4949 7590 4959 7642
rect 4959 7590 5005 7642
rect 4709 7588 4765 7590
rect 4789 7588 4845 7590
rect 4869 7588 4925 7590
rect 4949 7588 5005 7590
rect 4709 6554 4765 6556
rect 4789 6554 4845 6556
rect 4869 6554 4925 6556
rect 4949 6554 5005 6556
rect 4709 6502 4755 6554
rect 4755 6502 4765 6554
rect 4789 6502 4819 6554
rect 4819 6502 4831 6554
rect 4831 6502 4845 6554
rect 4869 6502 4883 6554
rect 4883 6502 4895 6554
rect 4895 6502 4925 6554
rect 4949 6502 4959 6554
rect 4959 6502 5005 6554
rect 4709 6500 4765 6502
rect 4789 6500 4845 6502
rect 4869 6500 4925 6502
rect 4949 6500 5005 6502
rect 4049 4922 4105 4924
rect 4129 4922 4185 4924
rect 4209 4922 4265 4924
rect 4289 4922 4345 4924
rect 4049 4870 4095 4922
rect 4095 4870 4105 4922
rect 4129 4870 4159 4922
rect 4159 4870 4171 4922
rect 4171 4870 4185 4922
rect 4209 4870 4223 4922
rect 4223 4870 4235 4922
rect 4235 4870 4265 4922
rect 4289 4870 4299 4922
rect 4299 4870 4345 4922
rect 4049 4868 4105 4870
rect 4129 4868 4185 4870
rect 4209 4868 4265 4870
rect 4289 4868 4345 4870
rect 4049 3834 4105 3836
rect 4129 3834 4185 3836
rect 4209 3834 4265 3836
rect 4289 3834 4345 3836
rect 4049 3782 4095 3834
rect 4095 3782 4105 3834
rect 4129 3782 4159 3834
rect 4159 3782 4171 3834
rect 4171 3782 4185 3834
rect 4209 3782 4223 3834
rect 4223 3782 4235 3834
rect 4235 3782 4265 3834
rect 4289 3782 4299 3834
rect 4299 3782 4345 3834
rect 4049 3780 4105 3782
rect 4129 3780 4185 3782
rect 4209 3780 4265 3782
rect 4289 3780 4345 3782
rect 4709 5466 4765 5468
rect 4789 5466 4845 5468
rect 4869 5466 4925 5468
rect 4949 5466 5005 5468
rect 4709 5414 4755 5466
rect 4755 5414 4765 5466
rect 4789 5414 4819 5466
rect 4819 5414 4831 5466
rect 4831 5414 4845 5466
rect 4869 5414 4883 5466
rect 4883 5414 4895 5466
rect 4895 5414 4925 5466
rect 4949 5414 4959 5466
rect 4959 5414 5005 5466
rect 4709 5412 4765 5414
rect 4789 5412 4845 5414
rect 4869 5412 4925 5414
rect 4949 5412 5005 5414
rect 4709 4378 4765 4380
rect 4789 4378 4845 4380
rect 4869 4378 4925 4380
rect 4949 4378 5005 4380
rect 4709 4326 4755 4378
rect 4755 4326 4765 4378
rect 4789 4326 4819 4378
rect 4819 4326 4831 4378
rect 4831 4326 4845 4378
rect 4869 4326 4883 4378
rect 4883 4326 4895 4378
rect 4895 4326 4925 4378
rect 4949 4326 4959 4378
rect 4959 4326 5005 4378
rect 4709 4324 4765 4326
rect 4789 4324 4845 4326
rect 4869 4324 4925 4326
rect 4949 4324 5005 4326
rect 4709 3290 4765 3292
rect 4789 3290 4845 3292
rect 4869 3290 4925 3292
rect 4949 3290 5005 3292
rect 4709 3238 4755 3290
rect 4755 3238 4765 3290
rect 4789 3238 4819 3290
rect 4819 3238 4831 3290
rect 4831 3238 4845 3290
rect 4869 3238 4883 3290
rect 4883 3238 4895 3290
rect 4895 3238 4925 3290
rect 4949 3238 4959 3290
rect 4959 3238 5005 3290
rect 4709 3236 4765 3238
rect 4789 3236 4845 3238
rect 4869 3236 4925 3238
rect 4949 3236 5005 3238
rect 2042 3052 2098 3088
rect 2042 3032 2044 3052
rect 2044 3032 2096 3052
rect 2096 3032 2098 3052
rect 1582 2080 1638 2136
rect 1306 1400 1362 1456
rect 4049 2746 4105 2748
rect 4129 2746 4185 2748
rect 4209 2746 4265 2748
rect 4289 2746 4345 2748
rect 4049 2694 4095 2746
rect 4095 2694 4105 2746
rect 4129 2694 4159 2746
rect 4159 2694 4171 2746
rect 4171 2694 4185 2746
rect 4209 2694 4223 2746
rect 4223 2694 4235 2746
rect 4235 2694 4265 2746
rect 4289 2694 4299 2746
rect 4299 2694 4345 2746
rect 4049 2692 4105 2694
rect 4129 2692 4185 2694
rect 4209 2692 4265 2694
rect 4289 2692 4345 2694
rect 5538 10512 5594 10568
rect 5354 6740 5356 6760
rect 5356 6740 5408 6760
rect 5408 6740 5410 6760
rect 5354 6704 5410 6740
rect 6090 12180 6092 12200
rect 6092 12180 6144 12200
rect 6144 12180 6146 12200
rect 6090 12144 6146 12180
rect 6458 13368 6514 13424
rect 6826 24812 6882 24848
rect 6826 24792 6828 24812
rect 6828 24792 6880 24812
rect 6880 24792 6882 24812
rect 6826 20168 6882 20224
rect 7286 19896 7342 19952
rect 5814 9560 5870 9616
rect 5722 6160 5778 6216
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 8574 25744 8630 25800
rect 7838 20712 7894 20768
rect 8758 23704 8814 23760
rect 7838 18672 7894 18728
rect 8482 20032 8538 20088
rect 10236 25594 10292 25596
rect 10316 25594 10372 25596
rect 10396 25594 10452 25596
rect 10476 25594 10532 25596
rect 10236 25542 10282 25594
rect 10282 25542 10292 25594
rect 10316 25542 10346 25594
rect 10346 25542 10358 25594
rect 10358 25542 10372 25594
rect 10396 25542 10410 25594
rect 10410 25542 10422 25594
rect 10422 25542 10452 25594
rect 10476 25542 10486 25594
rect 10486 25542 10532 25594
rect 10236 25540 10292 25542
rect 10316 25540 10372 25542
rect 10396 25540 10452 25542
rect 10476 25540 10532 25542
rect 10414 25356 10470 25392
rect 10414 25336 10416 25356
rect 10416 25336 10468 25356
rect 10468 25336 10470 25356
rect 9678 24656 9734 24712
rect 9770 23860 9826 23896
rect 9770 23840 9772 23860
rect 9772 23840 9824 23860
rect 9824 23840 9826 23860
rect 10236 24506 10292 24508
rect 10316 24506 10372 24508
rect 10396 24506 10452 24508
rect 10476 24506 10532 24508
rect 10236 24454 10282 24506
rect 10282 24454 10292 24506
rect 10316 24454 10346 24506
rect 10346 24454 10358 24506
rect 10358 24454 10372 24506
rect 10396 24454 10410 24506
rect 10410 24454 10422 24506
rect 10422 24454 10452 24506
rect 10476 24454 10486 24506
rect 10486 24454 10532 24506
rect 10236 24452 10292 24454
rect 10316 24452 10372 24454
rect 10396 24452 10452 24454
rect 10476 24452 10532 24454
rect 10506 23840 10562 23896
rect 10138 23704 10194 23760
rect 8850 20304 8906 20360
rect 9218 20168 9274 20224
rect 8298 19216 8354 19272
rect 8942 16532 8944 16552
rect 8944 16532 8996 16552
rect 8996 16532 8998 16552
rect 8942 16496 8998 16532
rect 9770 22752 9826 22808
rect 10236 23418 10292 23420
rect 10316 23418 10372 23420
rect 10396 23418 10452 23420
rect 10476 23418 10532 23420
rect 10236 23366 10282 23418
rect 10282 23366 10292 23418
rect 10316 23366 10346 23418
rect 10346 23366 10358 23418
rect 10358 23366 10372 23418
rect 10396 23366 10410 23418
rect 10410 23366 10422 23418
rect 10422 23366 10452 23418
rect 10476 23366 10486 23418
rect 10486 23366 10532 23418
rect 10236 23364 10292 23366
rect 10316 23364 10372 23366
rect 10396 23364 10452 23366
rect 10476 23364 10532 23366
rect 8850 15000 8906 15056
rect 8114 13232 8170 13288
rect 7654 7792 7710 7848
rect 7838 7112 7894 7168
rect 7930 6160 7986 6216
rect 3882 2372 3938 2408
rect 3882 2352 3884 2372
rect 3884 2352 3936 2372
rect 3936 2352 3938 2372
rect 4709 2202 4765 2204
rect 4789 2202 4845 2204
rect 4869 2202 4925 2204
rect 4949 2202 5005 2204
rect 4709 2150 4755 2202
rect 4755 2150 4765 2202
rect 4789 2150 4819 2202
rect 4819 2150 4831 2202
rect 4831 2150 4845 2202
rect 4869 2150 4883 2202
rect 4883 2150 4895 2202
rect 4895 2150 4925 2202
rect 4949 2150 4959 2202
rect 4959 2150 5005 2202
rect 4709 2148 4765 2150
rect 4789 2148 4845 2150
rect 4869 2148 4925 2150
rect 4949 2148 5005 2150
rect 9678 17740 9734 17776
rect 9678 17720 9680 17740
rect 9680 17720 9732 17740
rect 9732 17720 9734 17740
rect 9954 22072 10010 22128
rect 10236 22330 10292 22332
rect 10316 22330 10372 22332
rect 10396 22330 10452 22332
rect 10476 22330 10532 22332
rect 10236 22278 10282 22330
rect 10282 22278 10292 22330
rect 10316 22278 10346 22330
rect 10346 22278 10358 22330
rect 10358 22278 10372 22330
rect 10396 22278 10410 22330
rect 10410 22278 10422 22330
rect 10422 22278 10452 22330
rect 10476 22278 10486 22330
rect 10486 22278 10532 22330
rect 10236 22276 10292 22278
rect 10316 22276 10372 22278
rect 10396 22276 10452 22278
rect 10476 22276 10532 22278
rect 10230 22072 10286 22128
rect 10046 21528 10102 21584
rect 10236 21242 10292 21244
rect 10316 21242 10372 21244
rect 10396 21242 10452 21244
rect 10476 21242 10532 21244
rect 10236 21190 10282 21242
rect 10282 21190 10292 21242
rect 10316 21190 10346 21242
rect 10346 21190 10358 21242
rect 10358 21190 10372 21242
rect 10396 21190 10410 21242
rect 10410 21190 10422 21242
rect 10422 21190 10452 21242
rect 10476 21190 10486 21242
rect 10486 21190 10532 21242
rect 10236 21188 10292 21190
rect 10316 21188 10372 21190
rect 10396 21188 10452 21190
rect 10476 21188 10532 21190
rect 10236 20154 10292 20156
rect 10316 20154 10372 20156
rect 10396 20154 10452 20156
rect 10476 20154 10532 20156
rect 10236 20102 10282 20154
rect 10282 20102 10292 20154
rect 10316 20102 10346 20154
rect 10346 20102 10358 20154
rect 10358 20102 10372 20154
rect 10396 20102 10410 20154
rect 10410 20102 10422 20154
rect 10422 20102 10452 20154
rect 10476 20102 10486 20154
rect 10486 20102 10532 20154
rect 10236 20100 10292 20102
rect 10316 20100 10372 20102
rect 10396 20100 10452 20102
rect 10476 20100 10532 20102
rect 10896 26138 10952 26140
rect 10976 26138 11032 26140
rect 11056 26138 11112 26140
rect 11136 26138 11192 26140
rect 10896 26086 10942 26138
rect 10942 26086 10952 26138
rect 10976 26086 11006 26138
rect 11006 26086 11018 26138
rect 11018 26086 11032 26138
rect 11056 26086 11070 26138
rect 11070 26086 11082 26138
rect 11082 26086 11112 26138
rect 11136 26086 11146 26138
rect 11146 26086 11192 26138
rect 10896 26084 10952 26086
rect 10976 26084 11032 26086
rect 11056 26084 11112 26086
rect 11136 26084 11192 26086
rect 10896 25050 10952 25052
rect 10976 25050 11032 25052
rect 11056 25050 11112 25052
rect 11136 25050 11192 25052
rect 10896 24998 10942 25050
rect 10942 24998 10952 25050
rect 10976 24998 11006 25050
rect 11006 24998 11018 25050
rect 11018 24998 11032 25050
rect 11056 24998 11070 25050
rect 11070 24998 11082 25050
rect 11082 24998 11112 25050
rect 11136 24998 11146 25050
rect 11146 24998 11192 25050
rect 10896 24996 10952 24998
rect 10976 24996 11032 24998
rect 11056 24996 11112 24998
rect 11136 24996 11192 24998
rect 10896 23962 10952 23964
rect 10976 23962 11032 23964
rect 11056 23962 11112 23964
rect 11136 23962 11192 23964
rect 10896 23910 10942 23962
rect 10942 23910 10952 23962
rect 10976 23910 11006 23962
rect 11006 23910 11018 23962
rect 11018 23910 11032 23962
rect 11056 23910 11070 23962
rect 11070 23910 11082 23962
rect 11082 23910 11112 23962
rect 11136 23910 11146 23962
rect 11146 23910 11192 23962
rect 10896 23908 10952 23910
rect 10976 23908 11032 23910
rect 11056 23908 11112 23910
rect 11136 23908 11192 23910
rect 10896 22874 10952 22876
rect 10976 22874 11032 22876
rect 11056 22874 11112 22876
rect 11136 22874 11192 22876
rect 10896 22822 10942 22874
rect 10942 22822 10952 22874
rect 10976 22822 11006 22874
rect 11006 22822 11018 22874
rect 11018 22822 11032 22874
rect 11056 22822 11070 22874
rect 11070 22822 11082 22874
rect 11082 22822 11112 22874
rect 11136 22822 11146 22874
rect 11146 22822 11192 22874
rect 10896 22820 10952 22822
rect 10976 22820 11032 22822
rect 11056 22820 11112 22822
rect 11136 22820 11192 22822
rect 10782 21972 10784 21992
rect 10784 21972 10836 21992
rect 10836 21972 10838 21992
rect 10782 21936 10838 21972
rect 10896 21786 10952 21788
rect 10976 21786 11032 21788
rect 11056 21786 11112 21788
rect 11136 21786 11192 21788
rect 10896 21734 10942 21786
rect 10942 21734 10952 21786
rect 10976 21734 11006 21786
rect 11006 21734 11018 21786
rect 11018 21734 11032 21786
rect 11056 21734 11070 21786
rect 11070 21734 11082 21786
rect 11082 21734 11112 21786
rect 11136 21734 11146 21786
rect 11146 21734 11192 21786
rect 10896 21732 10952 21734
rect 10976 21732 11032 21734
rect 11056 21732 11112 21734
rect 11136 21732 11192 21734
rect 10690 20032 10746 20088
rect 10236 19066 10292 19068
rect 10316 19066 10372 19068
rect 10396 19066 10452 19068
rect 10476 19066 10532 19068
rect 10236 19014 10282 19066
rect 10282 19014 10292 19066
rect 10316 19014 10346 19066
rect 10346 19014 10358 19066
rect 10358 19014 10372 19066
rect 10396 19014 10410 19066
rect 10410 19014 10422 19066
rect 10422 19014 10452 19066
rect 10476 19014 10486 19066
rect 10486 19014 10532 19066
rect 10236 19012 10292 19014
rect 10316 19012 10372 19014
rect 10396 19012 10452 19014
rect 10476 19012 10532 19014
rect 10236 17978 10292 17980
rect 10316 17978 10372 17980
rect 10396 17978 10452 17980
rect 10476 17978 10532 17980
rect 10236 17926 10282 17978
rect 10282 17926 10292 17978
rect 10316 17926 10346 17978
rect 10346 17926 10358 17978
rect 10358 17926 10372 17978
rect 10396 17926 10410 17978
rect 10410 17926 10422 17978
rect 10422 17926 10452 17978
rect 10476 17926 10486 17978
rect 10486 17926 10532 17978
rect 10236 17924 10292 17926
rect 10316 17924 10372 17926
rect 10396 17924 10452 17926
rect 10476 17924 10532 17926
rect 10896 20698 10952 20700
rect 10976 20698 11032 20700
rect 11056 20698 11112 20700
rect 11136 20698 11192 20700
rect 10896 20646 10942 20698
rect 10942 20646 10952 20698
rect 10976 20646 11006 20698
rect 11006 20646 11018 20698
rect 11018 20646 11032 20698
rect 11056 20646 11070 20698
rect 11070 20646 11082 20698
rect 11082 20646 11112 20698
rect 11136 20646 11146 20698
rect 11146 20646 11192 20698
rect 10896 20644 10952 20646
rect 10976 20644 11032 20646
rect 11056 20644 11112 20646
rect 11136 20644 11192 20646
rect 11702 20304 11758 20360
rect 10896 19610 10952 19612
rect 10976 19610 11032 19612
rect 11056 19610 11112 19612
rect 11136 19610 11192 19612
rect 10896 19558 10942 19610
rect 10942 19558 10952 19610
rect 10976 19558 11006 19610
rect 11006 19558 11018 19610
rect 11018 19558 11032 19610
rect 11056 19558 11070 19610
rect 11070 19558 11082 19610
rect 11082 19558 11112 19610
rect 11136 19558 11146 19610
rect 11146 19558 11192 19610
rect 10896 19556 10952 19558
rect 10976 19556 11032 19558
rect 11056 19556 11112 19558
rect 11136 19556 11192 19558
rect 10966 18808 11022 18864
rect 10896 18522 10952 18524
rect 10976 18522 11032 18524
rect 11056 18522 11112 18524
rect 11136 18522 11192 18524
rect 10896 18470 10942 18522
rect 10942 18470 10952 18522
rect 10976 18470 11006 18522
rect 11006 18470 11018 18522
rect 11018 18470 11032 18522
rect 11056 18470 11070 18522
rect 11070 18470 11082 18522
rect 11082 18470 11112 18522
rect 11136 18470 11146 18522
rect 11146 18470 11192 18522
rect 10896 18468 10952 18470
rect 10976 18468 11032 18470
rect 11056 18468 11112 18470
rect 11136 18468 11192 18470
rect 9770 13232 9826 13288
rect 8206 7112 8262 7168
rect 9770 9424 9826 9480
rect 9678 9152 9734 9208
rect 9862 9016 9918 9072
rect 10236 16890 10292 16892
rect 10316 16890 10372 16892
rect 10396 16890 10452 16892
rect 10476 16890 10532 16892
rect 10236 16838 10282 16890
rect 10282 16838 10292 16890
rect 10316 16838 10346 16890
rect 10346 16838 10358 16890
rect 10358 16838 10372 16890
rect 10396 16838 10410 16890
rect 10410 16838 10422 16890
rect 10422 16838 10452 16890
rect 10476 16838 10486 16890
rect 10486 16838 10532 16890
rect 10236 16836 10292 16838
rect 10316 16836 10372 16838
rect 10396 16836 10452 16838
rect 10476 16836 10532 16838
rect 10506 16496 10562 16552
rect 10896 17434 10952 17436
rect 10976 17434 11032 17436
rect 11056 17434 11112 17436
rect 11136 17434 11192 17436
rect 10896 17382 10942 17434
rect 10942 17382 10952 17434
rect 10976 17382 11006 17434
rect 11006 17382 11018 17434
rect 11018 17382 11032 17434
rect 11056 17382 11070 17434
rect 11070 17382 11082 17434
rect 11082 17382 11112 17434
rect 11136 17382 11146 17434
rect 11146 17382 11192 17434
rect 10896 17380 10952 17382
rect 10976 17380 11032 17382
rect 11056 17380 11112 17382
rect 11136 17380 11192 17382
rect 10896 16346 10952 16348
rect 10976 16346 11032 16348
rect 11056 16346 11112 16348
rect 11136 16346 11192 16348
rect 10896 16294 10942 16346
rect 10942 16294 10952 16346
rect 10976 16294 11006 16346
rect 11006 16294 11018 16346
rect 11018 16294 11032 16346
rect 11056 16294 11070 16346
rect 11070 16294 11082 16346
rect 11082 16294 11112 16346
rect 11136 16294 11146 16346
rect 11146 16294 11192 16346
rect 10896 16292 10952 16294
rect 10976 16292 11032 16294
rect 11056 16292 11112 16294
rect 11136 16292 11192 16294
rect 10236 15802 10292 15804
rect 10316 15802 10372 15804
rect 10396 15802 10452 15804
rect 10476 15802 10532 15804
rect 10236 15750 10282 15802
rect 10282 15750 10292 15802
rect 10316 15750 10346 15802
rect 10346 15750 10358 15802
rect 10358 15750 10372 15802
rect 10396 15750 10410 15802
rect 10410 15750 10422 15802
rect 10422 15750 10452 15802
rect 10476 15750 10486 15802
rect 10486 15750 10532 15802
rect 10236 15748 10292 15750
rect 10316 15748 10372 15750
rect 10396 15748 10452 15750
rect 10476 15748 10532 15750
rect 10236 14714 10292 14716
rect 10316 14714 10372 14716
rect 10396 14714 10452 14716
rect 10476 14714 10532 14716
rect 10236 14662 10282 14714
rect 10282 14662 10292 14714
rect 10316 14662 10346 14714
rect 10346 14662 10358 14714
rect 10358 14662 10372 14714
rect 10396 14662 10410 14714
rect 10410 14662 10422 14714
rect 10422 14662 10452 14714
rect 10476 14662 10486 14714
rect 10486 14662 10532 14714
rect 10236 14660 10292 14662
rect 10316 14660 10372 14662
rect 10396 14660 10452 14662
rect 10476 14660 10532 14662
rect 10506 13776 10562 13832
rect 10236 13626 10292 13628
rect 10316 13626 10372 13628
rect 10396 13626 10452 13628
rect 10476 13626 10532 13628
rect 10236 13574 10282 13626
rect 10282 13574 10292 13626
rect 10316 13574 10346 13626
rect 10346 13574 10358 13626
rect 10358 13574 10372 13626
rect 10396 13574 10410 13626
rect 10410 13574 10422 13626
rect 10422 13574 10452 13626
rect 10476 13574 10486 13626
rect 10486 13574 10532 13626
rect 10236 13572 10292 13574
rect 10316 13572 10372 13574
rect 10396 13572 10452 13574
rect 10476 13572 10532 13574
rect 11426 16360 11482 16416
rect 11886 17584 11942 17640
rect 11242 15952 11298 16008
rect 12162 24248 12218 24304
rect 12346 19252 12348 19272
rect 12348 19252 12400 19272
rect 12400 19252 12402 19272
rect 12346 19216 12402 19252
rect 10896 15258 10952 15260
rect 10976 15258 11032 15260
rect 11056 15258 11112 15260
rect 11136 15258 11192 15260
rect 10896 15206 10942 15258
rect 10942 15206 10952 15258
rect 10976 15206 11006 15258
rect 11006 15206 11018 15258
rect 11018 15206 11032 15258
rect 11056 15206 11070 15258
rect 11070 15206 11082 15258
rect 11082 15206 11112 15258
rect 11136 15206 11146 15258
rect 11146 15206 11192 15258
rect 10896 15204 10952 15206
rect 10976 15204 11032 15206
rect 11056 15204 11112 15206
rect 11136 15204 11192 15206
rect 10896 14170 10952 14172
rect 10976 14170 11032 14172
rect 11056 14170 11112 14172
rect 11136 14170 11192 14172
rect 10896 14118 10942 14170
rect 10942 14118 10952 14170
rect 10976 14118 11006 14170
rect 11006 14118 11018 14170
rect 11018 14118 11032 14170
rect 11056 14118 11070 14170
rect 11070 14118 11082 14170
rect 11082 14118 11112 14170
rect 11136 14118 11146 14170
rect 11146 14118 11192 14170
rect 10896 14116 10952 14118
rect 10976 14116 11032 14118
rect 11056 14116 11112 14118
rect 11136 14116 11192 14118
rect 10782 13776 10838 13832
rect 10236 12538 10292 12540
rect 10316 12538 10372 12540
rect 10396 12538 10452 12540
rect 10476 12538 10532 12540
rect 10236 12486 10282 12538
rect 10282 12486 10292 12538
rect 10316 12486 10346 12538
rect 10346 12486 10358 12538
rect 10358 12486 10372 12538
rect 10396 12486 10410 12538
rect 10410 12486 10422 12538
rect 10422 12486 10452 12538
rect 10476 12486 10486 12538
rect 10486 12486 10532 12538
rect 10236 12484 10292 12486
rect 10316 12484 10372 12486
rect 10396 12484 10452 12486
rect 10476 12484 10532 12486
rect 10236 11450 10292 11452
rect 10316 11450 10372 11452
rect 10396 11450 10452 11452
rect 10476 11450 10532 11452
rect 10236 11398 10282 11450
rect 10282 11398 10292 11450
rect 10316 11398 10346 11450
rect 10346 11398 10358 11450
rect 10358 11398 10372 11450
rect 10396 11398 10410 11450
rect 10410 11398 10422 11450
rect 10422 11398 10452 11450
rect 10476 11398 10486 11450
rect 10486 11398 10532 11450
rect 10236 11396 10292 11398
rect 10316 11396 10372 11398
rect 10396 11396 10452 11398
rect 10476 11396 10532 11398
rect 10236 10362 10292 10364
rect 10316 10362 10372 10364
rect 10396 10362 10452 10364
rect 10476 10362 10532 10364
rect 10236 10310 10282 10362
rect 10282 10310 10292 10362
rect 10316 10310 10346 10362
rect 10346 10310 10358 10362
rect 10358 10310 10372 10362
rect 10396 10310 10410 10362
rect 10410 10310 10422 10362
rect 10422 10310 10452 10362
rect 10476 10310 10486 10362
rect 10486 10310 10532 10362
rect 10236 10308 10292 10310
rect 10316 10308 10372 10310
rect 10396 10308 10452 10310
rect 10476 10308 10532 10310
rect 10236 9274 10292 9276
rect 10316 9274 10372 9276
rect 10396 9274 10452 9276
rect 10476 9274 10532 9276
rect 10236 9222 10282 9274
rect 10282 9222 10292 9274
rect 10316 9222 10346 9274
rect 10346 9222 10358 9274
rect 10358 9222 10372 9274
rect 10396 9222 10410 9274
rect 10410 9222 10422 9274
rect 10422 9222 10452 9274
rect 10476 9222 10486 9274
rect 10486 9222 10532 9274
rect 10236 9220 10292 9222
rect 10316 9220 10372 9222
rect 10396 9220 10452 9222
rect 10476 9220 10532 9222
rect 9678 8880 9734 8936
rect 9586 6704 9642 6760
rect 9678 6316 9734 6352
rect 9678 6296 9680 6316
rect 9680 6296 9732 6316
rect 9732 6296 9734 6316
rect 9586 6160 9642 6216
rect 10138 9016 10194 9072
rect 9862 2896 9918 2952
rect 10236 8186 10292 8188
rect 10316 8186 10372 8188
rect 10396 8186 10452 8188
rect 10476 8186 10532 8188
rect 10236 8134 10282 8186
rect 10282 8134 10292 8186
rect 10316 8134 10346 8186
rect 10346 8134 10358 8186
rect 10358 8134 10372 8186
rect 10396 8134 10410 8186
rect 10410 8134 10422 8186
rect 10422 8134 10452 8186
rect 10476 8134 10486 8186
rect 10486 8134 10532 8186
rect 10236 8132 10292 8134
rect 10316 8132 10372 8134
rect 10396 8132 10452 8134
rect 10476 8132 10532 8134
rect 10236 7098 10292 7100
rect 10316 7098 10372 7100
rect 10396 7098 10452 7100
rect 10476 7098 10532 7100
rect 10236 7046 10282 7098
rect 10282 7046 10292 7098
rect 10316 7046 10346 7098
rect 10346 7046 10358 7098
rect 10358 7046 10372 7098
rect 10396 7046 10410 7098
rect 10410 7046 10422 7098
rect 10422 7046 10452 7098
rect 10476 7046 10486 7098
rect 10486 7046 10532 7098
rect 10236 7044 10292 7046
rect 10316 7044 10372 7046
rect 10396 7044 10452 7046
rect 10476 7044 10532 7046
rect 10236 6010 10292 6012
rect 10316 6010 10372 6012
rect 10396 6010 10452 6012
rect 10476 6010 10532 6012
rect 10236 5958 10282 6010
rect 10282 5958 10292 6010
rect 10316 5958 10346 6010
rect 10346 5958 10358 6010
rect 10358 5958 10372 6010
rect 10396 5958 10410 6010
rect 10410 5958 10422 6010
rect 10422 5958 10452 6010
rect 10476 5958 10486 6010
rect 10486 5958 10532 6010
rect 10236 5956 10292 5958
rect 10316 5956 10372 5958
rect 10396 5956 10452 5958
rect 10476 5956 10532 5958
rect 10236 4922 10292 4924
rect 10316 4922 10372 4924
rect 10396 4922 10452 4924
rect 10476 4922 10532 4924
rect 10236 4870 10282 4922
rect 10282 4870 10292 4922
rect 10316 4870 10346 4922
rect 10346 4870 10358 4922
rect 10358 4870 10372 4922
rect 10396 4870 10410 4922
rect 10410 4870 10422 4922
rect 10422 4870 10452 4922
rect 10476 4870 10486 4922
rect 10486 4870 10532 4922
rect 10236 4868 10292 4870
rect 10316 4868 10372 4870
rect 10396 4868 10452 4870
rect 10476 4868 10532 4870
rect 10236 3834 10292 3836
rect 10316 3834 10372 3836
rect 10396 3834 10452 3836
rect 10476 3834 10532 3836
rect 10236 3782 10282 3834
rect 10282 3782 10292 3834
rect 10316 3782 10346 3834
rect 10346 3782 10358 3834
rect 10358 3782 10372 3834
rect 10396 3782 10410 3834
rect 10410 3782 10422 3834
rect 10422 3782 10452 3834
rect 10476 3782 10486 3834
rect 10486 3782 10532 3834
rect 10236 3780 10292 3782
rect 10316 3780 10372 3782
rect 10396 3780 10452 3782
rect 10476 3780 10532 3782
rect 10236 2746 10292 2748
rect 10316 2746 10372 2748
rect 10396 2746 10452 2748
rect 10476 2746 10532 2748
rect 10236 2694 10282 2746
rect 10282 2694 10292 2746
rect 10316 2694 10346 2746
rect 10346 2694 10358 2746
rect 10358 2694 10372 2746
rect 10396 2694 10410 2746
rect 10410 2694 10422 2746
rect 10422 2694 10452 2746
rect 10476 2694 10486 2746
rect 10486 2694 10532 2746
rect 10236 2692 10292 2694
rect 10316 2692 10372 2694
rect 10396 2692 10452 2694
rect 10476 2692 10532 2694
rect 10896 13082 10952 13084
rect 10976 13082 11032 13084
rect 11056 13082 11112 13084
rect 11136 13082 11192 13084
rect 10896 13030 10942 13082
rect 10942 13030 10952 13082
rect 10976 13030 11006 13082
rect 11006 13030 11018 13082
rect 11018 13030 11032 13082
rect 11056 13030 11070 13082
rect 11070 13030 11082 13082
rect 11082 13030 11112 13082
rect 11136 13030 11146 13082
rect 11146 13030 11192 13082
rect 10896 13028 10952 13030
rect 10976 13028 11032 13030
rect 11056 13028 11112 13030
rect 11136 13028 11192 13030
rect 11518 13776 11574 13832
rect 11058 12280 11114 12336
rect 10896 11994 10952 11996
rect 10976 11994 11032 11996
rect 11056 11994 11112 11996
rect 11136 11994 11192 11996
rect 10896 11942 10942 11994
rect 10942 11942 10952 11994
rect 10976 11942 11006 11994
rect 11006 11942 11018 11994
rect 11018 11942 11032 11994
rect 11056 11942 11070 11994
rect 11070 11942 11082 11994
rect 11082 11942 11112 11994
rect 11136 11942 11146 11994
rect 11146 11942 11192 11994
rect 10896 11940 10952 11942
rect 10976 11940 11032 11942
rect 11056 11940 11112 11942
rect 11136 11940 11192 11942
rect 10896 10906 10952 10908
rect 10976 10906 11032 10908
rect 11056 10906 11112 10908
rect 11136 10906 11192 10908
rect 10896 10854 10942 10906
rect 10942 10854 10952 10906
rect 10976 10854 11006 10906
rect 11006 10854 11018 10906
rect 11018 10854 11032 10906
rect 11056 10854 11070 10906
rect 11070 10854 11082 10906
rect 11082 10854 11112 10906
rect 11136 10854 11146 10906
rect 11146 10854 11192 10906
rect 10896 10852 10952 10854
rect 10976 10852 11032 10854
rect 11056 10852 11112 10854
rect 11136 10852 11192 10854
rect 10896 9818 10952 9820
rect 10976 9818 11032 9820
rect 11056 9818 11112 9820
rect 11136 9818 11192 9820
rect 10896 9766 10942 9818
rect 10942 9766 10952 9818
rect 10976 9766 11006 9818
rect 11006 9766 11018 9818
rect 11018 9766 11032 9818
rect 11056 9766 11070 9818
rect 11070 9766 11082 9818
rect 11082 9766 11112 9818
rect 11136 9766 11146 9818
rect 11146 9766 11192 9818
rect 10896 9764 10952 9766
rect 10976 9764 11032 9766
rect 11056 9764 11112 9766
rect 11136 9764 11192 9766
rect 11058 9560 11114 9616
rect 10782 9288 10838 9344
rect 11242 9016 11298 9072
rect 10896 8730 10952 8732
rect 10976 8730 11032 8732
rect 11056 8730 11112 8732
rect 11136 8730 11192 8732
rect 10896 8678 10942 8730
rect 10942 8678 10952 8730
rect 10976 8678 11006 8730
rect 11006 8678 11018 8730
rect 11018 8678 11032 8730
rect 11056 8678 11070 8730
rect 11070 8678 11082 8730
rect 11082 8678 11112 8730
rect 11136 8678 11146 8730
rect 11146 8678 11192 8730
rect 10896 8676 10952 8678
rect 10976 8676 11032 8678
rect 11056 8676 11112 8678
rect 11136 8676 11192 8678
rect 10896 7642 10952 7644
rect 10976 7642 11032 7644
rect 11056 7642 11112 7644
rect 11136 7642 11192 7644
rect 10896 7590 10942 7642
rect 10942 7590 10952 7642
rect 10976 7590 11006 7642
rect 11006 7590 11018 7642
rect 11018 7590 11032 7642
rect 11056 7590 11070 7642
rect 11070 7590 11082 7642
rect 11082 7590 11112 7642
rect 11136 7590 11146 7642
rect 11146 7590 11192 7642
rect 10896 7588 10952 7590
rect 10976 7588 11032 7590
rect 11056 7588 11112 7590
rect 11136 7588 11192 7590
rect 10896 6554 10952 6556
rect 10976 6554 11032 6556
rect 11056 6554 11112 6556
rect 11136 6554 11192 6556
rect 10896 6502 10942 6554
rect 10942 6502 10952 6554
rect 10976 6502 11006 6554
rect 11006 6502 11018 6554
rect 11018 6502 11032 6554
rect 11056 6502 11070 6554
rect 11070 6502 11082 6554
rect 11082 6502 11112 6554
rect 11136 6502 11146 6554
rect 11146 6502 11192 6554
rect 10896 6500 10952 6502
rect 10976 6500 11032 6502
rect 11056 6500 11112 6502
rect 11136 6500 11192 6502
rect 10896 5466 10952 5468
rect 10976 5466 11032 5468
rect 11056 5466 11112 5468
rect 11136 5466 11192 5468
rect 10896 5414 10942 5466
rect 10942 5414 10952 5466
rect 10976 5414 11006 5466
rect 11006 5414 11018 5466
rect 11018 5414 11032 5466
rect 11056 5414 11070 5466
rect 11070 5414 11082 5466
rect 11082 5414 11112 5466
rect 11136 5414 11146 5466
rect 11146 5414 11192 5466
rect 10896 5412 10952 5414
rect 10976 5412 11032 5414
rect 11056 5412 11112 5414
rect 11136 5412 11192 5414
rect 10896 4378 10952 4380
rect 10976 4378 11032 4380
rect 11056 4378 11112 4380
rect 11136 4378 11192 4380
rect 10896 4326 10942 4378
rect 10942 4326 10952 4378
rect 10976 4326 11006 4378
rect 11006 4326 11018 4378
rect 11018 4326 11032 4378
rect 11056 4326 11070 4378
rect 11070 4326 11082 4378
rect 11082 4326 11112 4378
rect 11136 4326 11146 4378
rect 11146 4326 11192 4378
rect 10896 4324 10952 4326
rect 10976 4324 11032 4326
rect 11056 4324 11112 4326
rect 11136 4324 11192 4326
rect 10896 3290 10952 3292
rect 10976 3290 11032 3292
rect 11056 3290 11112 3292
rect 11136 3290 11192 3292
rect 10896 3238 10942 3290
rect 10942 3238 10952 3290
rect 10976 3238 11006 3290
rect 11006 3238 11018 3290
rect 11018 3238 11032 3290
rect 11056 3238 11070 3290
rect 11070 3238 11082 3290
rect 11082 3238 11112 3290
rect 11136 3238 11146 3290
rect 11146 3238 11192 3290
rect 10896 3236 10952 3238
rect 10976 3236 11032 3238
rect 11056 3236 11112 3238
rect 11136 3236 11192 3238
rect 11886 12844 11942 12880
rect 11886 12824 11888 12844
rect 11888 12824 11940 12844
rect 11940 12824 11942 12844
rect 11886 12280 11942 12336
rect 12070 13812 12072 13832
rect 12072 13812 12124 13832
rect 12124 13812 12126 13832
rect 12070 13776 12126 13812
rect 12622 19252 12624 19272
rect 12624 19252 12676 19272
rect 12676 19252 12678 19272
rect 12622 19216 12678 19252
rect 12530 16496 12586 16552
rect 11978 12144 12034 12200
rect 11610 9424 11666 9480
rect 12714 12688 12770 12744
rect 16423 26682 16479 26684
rect 16503 26682 16559 26684
rect 16583 26682 16639 26684
rect 16663 26682 16719 26684
rect 16423 26630 16469 26682
rect 16469 26630 16479 26682
rect 16503 26630 16533 26682
rect 16533 26630 16545 26682
rect 16545 26630 16559 26682
rect 16583 26630 16597 26682
rect 16597 26630 16609 26682
rect 16609 26630 16639 26682
rect 16663 26630 16673 26682
rect 16673 26630 16719 26682
rect 16423 26628 16479 26630
rect 16503 26628 16559 26630
rect 16583 26628 16639 26630
rect 16663 26628 16719 26630
rect 14370 24112 14426 24168
rect 12990 20032 13046 20088
rect 11886 9152 11942 9208
rect 11886 8744 11942 8800
rect 12254 8744 12310 8800
rect 12530 9832 12586 9888
rect 12530 9696 12586 9752
rect 12898 10240 12954 10296
rect 12622 9424 12678 9480
rect 10896 2202 10952 2204
rect 10976 2202 11032 2204
rect 11056 2202 11112 2204
rect 11136 2202 11192 2204
rect 10896 2150 10942 2202
rect 10942 2150 10952 2202
rect 10976 2150 11006 2202
rect 11006 2150 11018 2202
rect 11018 2150 11032 2202
rect 11056 2150 11070 2202
rect 11070 2150 11082 2202
rect 11082 2150 11112 2202
rect 11136 2150 11146 2202
rect 11146 2150 11192 2202
rect 10896 2148 10952 2150
rect 10976 2148 11032 2150
rect 11056 2148 11112 2150
rect 11136 2148 11192 2150
rect 12806 2896 12862 2952
rect 13818 16632 13874 16688
rect 14554 23704 14610 23760
rect 14002 14320 14058 14376
rect 14646 18944 14702 19000
rect 14738 18692 14794 18728
rect 14738 18672 14740 18692
rect 14740 18672 14792 18692
rect 14792 18672 14794 18692
rect 15842 25744 15898 25800
rect 16423 25594 16479 25596
rect 16503 25594 16559 25596
rect 16583 25594 16639 25596
rect 16663 25594 16719 25596
rect 16423 25542 16469 25594
rect 16469 25542 16479 25594
rect 16503 25542 16533 25594
rect 16533 25542 16545 25594
rect 16545 25542 16559 25594
rect 16583 25542 16597 25594
rect 16597 25542 16609 25594
rect 16609 25542 16639 25594
rect 16663 25542 16673 25594
rect 16673 25542 16719 25594
rect 16423 25540 16479 25542
rect 16503 25540 16559 25542
rect 16583 25540 16639 25542
rect 16663 25540 16719 25542
rect 17083 26138 17139 26140
rect 17163 26138 17219 26140
rect 17243 26138 17299 26140
rect 17323 26138 17379 26140
rect 17083 26086 17129 26138
rect 17129 26086 17139 26138
rect 17163 26086 17193 26138
rect 17193 26086 17205 26138
rect 17205 26086 17219 26138
rect 17243 26086 17257 26138
rect 17257 26086 17269 26138
rect 17269 26086 17299 26138
rect 17323 26086 17333 26138
rect 17333 26086 17379 26138
rect 17083 26084 17139 26086
rect 17163 26084 17219 26086
rect 17243 26084 17299 26086
rect 17323 26084 17379 26086
rect 16423 24506 16479 24508
rect 16503 24506 16559 24508
rect 16583 24506 16639 24508
rect 16663 24506 16719 24508
rect 16423 24454 16469 24506
rect 16469 24454 16479 24506
rect 16503 24454 16533 24506
rect 16533 24454 16545 24506
rect 16545 24454 16559 24506
rect 16583 24454 16597 24506
rect 16597 24454 16609 24506
rect 16609 24454 16639 24506
rect 16663 24454 16673 24506
rect 16673 24454 16719 24506
rect 16423 24452 16479 24454
rect 16503 24452 16559 24454
rect 16583 24452 16639 24454
rect 16663 24452 16719 24454
rect 16394 24248 16450 24304
rect 15198 21528 15254 21584
rect 15106 19916 15162 19952
rect 15106 19896 15108 19916
rect 15108 19896 15160 19916
rect 15160 19896 15162 19916
rect 16423 23418 16479 23420
rect 16503 23418 16559 23420
rect 16583 23418 16639 23420
rect 16663 23418 16719 23420
rect 16423 23366 16469 23418
rect 16469 23366 16479 23418
rect 16503 23366 16533 23418
rect 16533 23366 16545 23418
rect 16545 23366 16559 23418
rect 16583 23366 16597 23418
rect 16597 23366 16609 23418
rect 16609 23366 16639 23418
rect 16663 23366 16673 23418
rect 16673 23366 16719 23418
rect 16423 23364 16479 23366
rect 16503 23364 16559 23366
rect 16583 23364 16639 23366
rect 16663 23364 16719 23366
rect 16423 22330 16479 22332
rect 16503 22330 16559 22332
rect 16583 22330 16639 22332
rect 16663 22330 16719 22332
rect 16423 22278 16469 22330
rect 16469 22278 16479 22330
rect 16503 22278 16533 22330
rect 16533 22278 16545 22330
rect 16545 22278 16559 22330
rect 16583 22278 16597 22330
rect 16597 22278 16609 22330
rect 16609 22278 16639 22330
rect 16663 22278 16673 22330
rect 16673 22278 16719 22330
rect 16423 22276 16479 22278
rect 16503 22276 16559 22278
rect 16583 22276 16639 22278
rect 16663 22276 16719 22278
rect 17083 25050 17139 25052
rect 17163 25050 17219 25052
rect 17243 25050 17299 25052
rect 17323 25050 17379 25052
rect 17083 24998 17129 25050
rect 17129 24998 17139 25050
rect 17163 24998 17193 25050
rect 17193 24998 17205 25050
rect 17205 24998 17219 25050
rect 17243 24998 17257 25050
rect 17257 24998 17269 25050
rect 17269 24998 17299 25050
rect 17323 24998 17333 25050
rect 17333 24998 17379 25050
rect 17083 24996 17139 24998
rect 17163 24996 17219 24998
rect 17243 24996 17299 24998
rect 17323 24996 17379 24998
rect 17498 24148 17500 24168
rect 17500 24148 17552 24168
rect 17552 24148 17554 24168
rect 17498 24112 17554 24148
rect 17083 23962 17139 23964
rect 17163 23962 17219 23964
rect 17243 23962 17299 23964
rect 17323 23962 17379 23964
rect 17083 23910 17129 23962
rect 17129 23910 17139 23962
rect 17163 23910 17193 23962
rect 17193 23910 17205 23962
rect 17205 23910 17219 23962
rect 17243 23910 17257 23962
rect 17257 23910 17269 23962
rect 17269 23910 17299 23962
rect 17323 23910 17333 23962
rect 17333 23910 17379 23962
rect 17083 23908 17139 23910
rect 17163 23908 17219 23910
rect 17243 23908 17299 23910
rect 17323 23908 17379 23910
rect 17083 22874 17139 22876
rect 17163 22874 17219 22876
rect 17243 22874 17299 22876
rect 17323 22874 17379 22876
rect 17083 22822 17129 22874
rect 17129 22822 17139 22874
rect 17163 22822 17193 22874
rect 17193 22822 17205 22874
rect 17205 22822 17219 22874
rect 17243 22822 17257 22874
rect 17257 22822 17269 22874
rect 17269 22822 17299 22874
rect 17323 22822 17333 22874
rect 17333 22822 17379 22874
rect 17083 22820 17139 22822
rect 17163 22820 17219 22822
rect 17243 22820 17299 22822
rect 17323 22820 17379 22822
rect 17590 22072 17646 22128
rect 16423 21242 16479 21244
rect 16503 21242 16559 21244
rect 16583 21242 16639 21244
rect 16663 21242 16719 21244
rect 16423 21190 16469 21242
rect 16469 21190 16479 21242
rect 16503 21190 16533 21242
rect 16533 21190 16545 21242
rect 16545 21190 16559 21242
rect 16583 21190 16597 21242
rect 16597 21190 16609 21242
rect 16609 21190 16639 21242
rect 16663 21190 16673 21242
rect 16673 21190 16719 21242
rect 16423 21188 16479 21190
rect 16503 21188 16559 21190
rect 16583 21188 16639 21190
rect 16663 21188 16719 21190
rect 15106 18284 15162 18320
rect 15106 18264 15108 18284
rect 15108 18264 15160 18284
rect 15160 18264 15162 18284
rect 15842 18964 15898 19000
rect 15842 18944 15844 18964
rect 15844 18944 15896 18964
rect 15896 18944 15898 18964
rect 15658 18672 15714 18728
rect 16423 20154 16479 20156
rect 16503 20154 16559 20156
rect 16583 20154 16639 20156
rect 16663 20154 16719 20156
rect 16423 20102 16469 20154
rect 16469 20102 16479 20154
rect 16503 20102 16533 20154
rect 16533 20102 16545 20154
rect 16545 20102 16559 20154
rect 16583 20102 16597 20154
rect 16597 20102 16609 20154
rect 16609 20102 16639 20154
rect 16663 20102 16673 20154
rect 16673 20102 16719 20154
rect 16423 20100 16479 20102
rect 16503 20100 16559 20102
rect 16583 20100 16639 20102
rect 16663 20100 16719 20102
rect 16423 19066 16479 19068
rect 16503 19066 16559 19068
rect 16583 19066 16639 19068
rect 16663 19066 16719 19068
rect 16423 19014 16469 19066
rect 16469 19014 16479 19066
rect 16503 19014 16533 19066
rect 16533 19014 16545 19066
rect 16545 19014 16559 19066
rect 16583 19014 16597 19066
rect 16597 19014 16609 19066
rect 16609 19014 16639 19066
rect 16663 19014 16673 19066
rect 16673 19014 16719 19066
rect 16423 19012 16479 19014
rect 16503 19012 16559 19014
rect 16583 19012 16639 19014
rect 16663 19012 16719 19014
rect 16670 18264 16726 18320
rect 17083 21786 17139 21788
rect 17163 21786 17219 21788
rect 17243 21786 17299 21788
rect 17323 21786 17379 21788
rect 17083 21734 17129 21786
rect 17129 21734 17139 21786
rect 17163 21734 17193 21786
rect 17193 21734 17205 21786
rect 17205 21734 17219 21786
rect 17243 21734 17257 21786
rect 17257 21734 17269 21786
rect 17269 21734 17299 21786
rect 17323 21734 17333 21786
rect 17333 21734 17379 21786
rect 17083 21732 17139 21734
rect 17163 21732 17219 21734
rect 17243 21732 17299 21734
rect 17323 21732 17379 21734
rect 17083 20698 17139 20700
rect 17163 20698 17219 20700
rect 17243 20698 17299 20700
rect 17323 20698 17379 20700
rect 17083 20646 17129 20698
rect 17129 20646 17139 20698
rect 17163 20646 17193 20698
rect 17193 20646 17205 20698
rect 17205 20646 17219 20698
rect 17243 20646 17257 20698
rect 17257 20646 17269 20698
rect 17269 20646 17299 20698
rect 17323 20646 17333 20698
rect 17333 20646 17379 20698
rect 17083 20644 17139 20646
rect 17163 20644 17219 20646
rect 17243 20644 17299 20646
rect 17323 20644 17379 20646
rect 17866 21936 17922 21992
rect 17083 19610 17139 19612
rect 17163 19610 17219 19612
rect 17243 19610 17299 19612
rect 17323 19610 17379 19612
rect 17083 19558 17129 19610
rect 17129 19558 17139 19610
rect 17163 19558 17193 19610
rect 17193 19558 17205 19610
rect 17205 19558 17219 19610
rect 17243 19558 17257 19610
rect 17257 19558 17269 19610
rect 17269 19558 17299 19610
rect 17323 19558 17333 19610
rect 17333 19558 17379 19610
rect 17083 19556 17139 19558
rect 17163 19556 17219 19558
rect 17243 19556 17299 19558
rect 17323 19556 17379 19558
rect 17083 18522 17139 18524
rect 17163 18522 17219 18524
rect 17243 18522 17299 18524
rect 17323 18522 17379 18524
rect 17083 18470 17129 18522
rect 17129 18470 17139 18522
rect 17163 18470 17193 18522
rect 17193 18470 17205 18522
rect 17205 18470 17219 18522
rect 17243 18470 17257 18522
rect 17257 18470 17269 18522
rect 17269 18470 17299 18522
rect 17323 18470 17333 18522
rect 17333 18470 17379 18522
rect 17083 18468 17139 18470
rect 17163 18468 17219 18470
rect 17243 18468 17299 18470
rect 17323 18468 17379 18470
rect 16423 17978 16479 17980
rect 16503 17978 16559 17980
rect 16583 17978 16639 17980
rect 16663 17978 16719 17980
rect 16423 17926 16469 17978
rect 16469 17926 16479 17978
rect 16503 17926 16533 17978
rect 16533 17926 16545 17978
rect 16545 17926 16559 17978
rect 16583 17926 16597 17978
rect 16597 17926 16609 17978
rect 16609 17926 16639 17978
rect 16663 17926 16673 17978
rect 16673 17926 16719 17978
rect 16423 17924 16479 17926
rect 16503 17924 16559 17926
rect 16583 17924 16639 17926
rect 16663 17924 16719 17926
rect 15198 15036 15200 15056
rect 15200 15036 15252 15056
rect 15252 15036 15254 15056
rect 15198 15000 15254 15036
rect 13910 11056 13966 11112
rect 13266 9696 13322 9752
rect 13174 9560 13230 9616
rect 13450 9424 13506 9480
rect 13542 9152 13598 9208
rect 13542 9016 13598 9072
rect 14830 10240 14886 10296
rect 14278 9288 14334 9344
rect 16423 16890 16479 16892
rect 16503 16890 16559 16892
rect 16583 16890 16639 16892
rect 16663 16890 16719 16892
rect 16423 16838 16469 16890
rect 16469 16838 16479 16890
rect 16503 16838 16533 16890
rect 16533 16838 16545 16890
rect 16545 16838 16559 16890
rect 16583 16838 16597 16890
rect 16597 16838 16609 16890
rect 16609 16838 16639 16890
rect 16663 16838 16673 16890
rect 16673 16838 16719 16890
rect 16423 16836 16479 16838
rect 16503 16836 16559 16838
rect 16583 16836 16639 16838
rect 16663 16836 16719 16838
rect 16423 15802 16479 15804
rect 16503 15802 16559 15804
rect 16583 15802 16639 15804
rect 16663 15802 16719 15804
rect 16423 15750 16469 15802
rect 16469 15750 16479 15802
rect 16503 15750 16533 15802
rect 16533 15750 16545 15802
rect 16545 15750 16559 15802
rect 16583 15750 16597 15802
rect 16597 15750 16609 15802
rect 16609 15750 16639 15802
rect 16663 15750 16673 15802
rect 16673 15750 16719 15802
rect 16423 15748 16479 15750
rect 16503 15748 16559 15750
rect 16583 15748 16639 15750
rect 16663 15748 16719 15750
rect 15842 12688 15898 12744
rect 15842 11600 15898 11656
rect 14462 5228 14518 5264
rect 14462 5208 14464 5228
rect 14464 5208 14516 5228
rect 14516 5208 14518 5228
rect 16423 14714 16479 14716
rect 16503 14714 16559 14716
rect 16583 14714 16639 14716
rect 16663 14714 16719 14716
rect 16423 14662 16469 14714
rect 16469 14662 16479 14714
rect 16503 14662 16533 14714
rect 16533 14662 16545 14714
rect 16545 14662 16559 14714
rect 16583 14662 16597 14714
rect 16597 14662 16609 14714
rect 16609 14662 16639 14714
rect 16663 14662 16673 14714
rect 16673 14662 16719 14714
rect 16423 14660 16479 14662
rect 16503 14660 16559 14662
rect 16583 14660 16639 14662
rect 16663 14660 16719 14662
rect 17083 17434 17139 17436
rect 17163 17434 17219 17436
rect 17243 17434 17299 17436
rect 17323 17434 17379 17436
rect 17083 17382 17129 17434
rect 17129 17382 17139 17434
rect 17163 17382 17193 17434
rect 17193 17382 17205 17434
rect 17205 17382 17219 17434
rect 17243 17382 17257 17434
rect 17257 17382 17269 17434
rect 17269 17382 17299 17434
rect 17323 17382 17333 17434
rect 17333 17382 17379 17434
rect 17083 17380 17139 17382
rect 17163 17380 17219 17382
rect 17243 17380 17299 17382
rect 17323 17380 17379 17382
rect 17083 16346 17139 16348
rect 17163 16346 17219 16348
rect 17243 16346 17299 16348
rect 17323 16346 17379 16348
rect 17083 16294 17129 16346
rect 17129 16294 17139 16346
rect 17163 16294 17193 16346
rect 17193 16294 17205 16346
rect 17205 16294 17219 16346
rect 17243 16294 17257 16346
rect 17257 16294 17269 16346
rect 17269 16294 17299 16346
rect 17323 16294 17333 16346
rect 17333 16294 17379 16346
rect 17083 16292 17139 16294
rect 17163 16292 17219 16294
rect 17243 16292 17299 16294
rect 17323 16292 17379 16294
rect 17083 15258 17139 15260
rect 17163 15258 17219 15260
rect 17243 15258 17299 15260
rect 17323 15258 17379 15260
rect 17083 15206 17129 15258
rect 17129 15206 17139 15258
rect 17163 15206 17193 15258
rect 17193 15206 17205 15258
rect 17205 15206 17219 15258
rect 17243 15206 17257 15258
rect 17257 15206 17269 15258
rect 17269 15206 17299 15258
rect 17323 15206 17333 15258
rect 17333 15206 17379 15258
rect 17083 15204 17139 15206
rect 17163 15204 17219 15206
rect 17243 15204 17299 15206
rect 17323 15204 17379 15206
rect 17083 14170 17139 14172
rect 17163 14170 17219 14172
rect 17243 14170 17299 14172
rect 17323 14170 17379 14172
rect 17083 14118 17129 14170
rect 17129 14118 17139 14170
rect 17163 14118 17193 14170
rect 17193 14118 17205 14170
rect 17205 14118 17219 14170
rect 17243 14118 17257 14170
rect 17257 14118 17269 14170
rect 17269 14118 17299 14170
rect 17323 14118 17333 14170
rect 17333 14118 17379 14170
rect 17083 14116 17139 14118
rect 17163 14116 17219 14118
rect 17243 14116 17299 14118
rect 17323 14116 17379 14118
rect 16423 13626 16479 13628
rect 16503 13626 16559 13628
rect 16583 13626 16639 13628
rect 16663 13626 16719 13628
rect 16423 13574 16469 13626
rect 16469 13574 16479 13626
rect 16503 13574 16533 13626
rect 16533 13574 16545 13626
rect 16545 13574 16559 13626
rect 16583 13574 16597 13626
rect 16597 13574 16609 13626
rect 16609 13574 16639 13626
rect 16663 13574 16673 13626
rect 16673 13574 16719 13626
rect 16423 13572 16479 13574
rect 16503 13572 16559 13574
rect 16583 13572 16639 13574
rect 16663 13572 16719 13574
rect 16578 13368 16634 13424
rect 17083 13082 17139 13084
rect 17163 13082 17219 13084
rect 17243 13082 17299 13084
rect 17323 13082 17379 13084
rect 17083 13030 17129 13082
rect 17129 13030 17139 13082
rect 17163 13030 17193 13082
rect 17193 13030 17205 13082
rect 17205 13030 17219 13082
rect 17243 13030 17257 13082
rect 17257 13030 17269 13082
rect 17269 13030 17299 13082
rect 17323 13030 17333 13082
rect 17333 13030 17379 13082
rect 17083 13028 17139 13030
rect 17163 13028 17219 13030
rect 17243 13028 17299 13030
rect 17323 13028 17379 13030
rect 16423 12538 16479 12540
rect 16503 12538 16559 12540
rect 16583 12538 16639 12540
rect 16663 12538 16719 12540
rect 16423 12486 16469 12538
rect 16469 12486 16479 12538
rect 16503 12486 16533 12538
rect 16533 12486 16545 12538
rect 16545 12486 16559 12538
rect 16583 12486 16597 12538
rect 16597 12486 16609 12538
rect 16609 12486 16639 12538
rect 16663 12486 16673 12538
rect 16673 12486 16719 12538
rect 16423 12484 16479 12486
rect 16503 12484 16559 12486
rect 16583 12484 16639 12486
rect 16663 12484 16719 12486
rect 16423 11450 16479 11452
rect 16503 11450 16559 11452
rect 16583 11450 16639 11452
rect 16663 11450 16719 11452
rect 16423 11398 16469 11450
rect 16469 11398 16479 11450
rect 16503 11398 16533 11450
rect 16533 11398 16545 11450
rect 16545 11398 16559 11450
rect 16583 11398 16597 11450
rect 16597 11398 16609 11450
rect 16609 11398 16639 11450
rect 16663 11398 16673 11450
rect 16673 11398 16719 11450
rect 16423 11396 16479 11398
rect 16503 11396 16559 11398
rect 16583 11396 16639 11398
rect 16663 11396 16719 11398
rect 16423 10362 16479 10364
rect 16503 10362 16559 10364
rect 16583 10362 16639 10364
rect 16663 10362 16719 10364
rect 16423 10310 16469 10362
rect 16469 10310 16479 10362
rect 16503 10310 16533 10362
rect 16533 10310 16545 10362
rect 16545 10310 16559 10362
rect 16583 10310 16597 10362
rect 16597 10310 16609 10362
rect 16609 10310 16639 10362
rect 16663 10310 16673 10362
rect 16673 10310 16719 10362
rect 16423 10308 16479 10310
rect 16503 10308 16559 10310
rect 16583 10308 16639 10310
rect 16663 10308 16719 10310
rect 16394 9696 16450 9752
rect 16578 9832 16634 9888
rect 16670 9696 16726 9752
rect 22926 28600 22982 28656
rect 18510 25356 18566 25392
rect 18510 25336 18512 25356
rect 18512 25336 18564 25356
rect 18564 25336 18566 25356
rect 22610 26682 22666 26684
rect 22690 26682 22746 26684
rect 22770 26682 22826 26684
rect 22850 26682 22906 26684
rect 22610 26630 22656 26682
rect 22656 26630 22666 26682
rect 22690 26630 22720 26682
rect 22720 26630 22732 26682
rect 22732 26630 22746 26682
rect 22770 26630 22784 26682
rect 22784 26630 22796 26682
rect 22796 26630 22826 26682
rect 22850 26630 22860 26682
rect 22860 26630 22906 26682
rect 22610 26628 22666 26630
rect 22690 26628 22746 26630
rect 22770 26628 22826 26630
rect 22850 26628 22906 26630
rect 18878 20304 18934 20360
rect 18418 16532 18420 16552
rect 18420 16532 18472 16552
rect 18472 16532 18474 16552
rect 18418 16496 18474 16532
rect 17083 11994 17139 11996
rect 17163 11994 17219 11996
rect 17243 11994 17299 11996
rect 17323 11994 17379 11996
rect 17083 11942 17129 11994
rect 17129 11942 17139 11994
rect 17163 11942 17193 11994
rect 17193 11942 17205 11994
rect 17205 11942 17219 11994
rect 17243 11942 17257 11994
rect 17257 11942 17269 11994
rect 17269 11942 17299 11994
rect 17323 11942 17333 11994
rect 17333 11942 17379 11994
rect 17083 11940 17139 11942
rect 17163 11940 17219 11942
rect 17243 11940 17299 11942
rect 17323 11940 17379 11942
rect 17314 11076 17370 11112
rect 17314 11056 17316 11076
rect 17316 11056 17368 11076
rect 17368 11056 17370 11076
rect 17083 10906 17139 10908
rect 17163 10906 17219 10908
rect 17243 10906 17299 10908
rect 17323 10906 17379 10908
rect 17083 10854 17129 10906
rect 17129 10854 17139 10906
rect 17163 10854 17193 10906
rect 17193 10854 17205 10906
rect 17205 10854 17219 10906
rect 17243 10854 17257 10906
rect 17257 10854 17269 10906
rect 17269 10854 17299 10906
rect 17323 10854 17333 10906
rect 17333 10854 17379 10906
rect 17083 10852 17139 10854
rect 17163 10852 17219 10854
rect 17243 10852 17299 10854
rect 17323 10852 17379 10854
rect 17130 10512 17186 10568
rect 18786 19216 18842 19272
rect 19430 19352 19486 19408
rect 21086 24792 21142 24848
rect 21270 23568 21326 23624
rect 18970 17992 19026 18048
rect 18970 16632 19026 16688
rect 19614 17040 19670 17096
rect 16946 9832 17002 9888
rect 17083 9818 17139 9820
rect 17163 9818 17219 9820
rect 17243 9818 17299 9820
rect 17323 9818 17379 9820
rect 17083 9766 17129 9818
rect 17129 9766 17139 9818
rect 17163 9766 17193 9818
rect 17193 9766 17205 9818
rect 17205 9766 17219 9818
rect 17243 9766 17257 9818
rect 17257 9766 17269 9818
rect 17269 9766 17299 9818
rect 17323 9766 17333 9818
rect 17333 9766 17379 9818
rect 17083 9764 17139 9766
rect 17163 9764 17219 9766
rect 17243 9764 17299 9766
rect 17323 9764 17379 9766
rect 16423 9274 16479 9276
rect 16503 9274 16559 9276
rect 16583 9274 16639 9276
rect 16663 9274 16719 9276
rect 16423 9222 16469 9274
rect 16469 9222 16479 9274
rect 16503 9222 16533 9274
rect 16533 9222 16545 9274
rect 16545 9222 16559 9274
rect 16583 9222 16597 9274
rect 16597 9222 16609 9274
rect 16609 9222 16639 9274
rect 16663 9222 16673 9274
rect 16673 9222 16719 9274
rect 16423 9220 16479 9222
rect 16503 9220 16559 9222
rect 16583 9220 16639 9222
rect 16663 9220 16719 9222
rect 16423 8186 16479 8188
rect 16503 8186 16559 8188
rect 16583 8186 16639 8188
rect 16663 8186 16719 8188
rect 16423 8134 16469 8186
rect 16469 8134 16479 8186
rect 16503 8134 16533 8186
rect 16533 8134 16545 8186
rect 16545 8134 16559 8186
rect 16583 8134 16597 8186
rect 16597 8134 16609 8186
rect 16609 8134 16639 8186
rect 16663 8134 16673 8186
rect 16673 8134 16719 8186
rect 16423 8132 16479 8134
rect 16503 8132 16559 8134
rect 16583 8132 16639 8134
rect 16663 8132 16719 8134
rect 15750 6296 15806 6352
rect 15566 4664 15622 4720
rect 15198 2624 15254 2680
rect 16423 7098 16479 7100
rect 16503 7098 16559 7100
rect 16583 7098 16639 7100
rect 16663 7098 16719 7100
rect 16423 7046 16469 7098
rect 16469 7046 16479 7098
rect 16503 7046 16533 7098
rect 16533 7046 16545 7098
rect 16545 7046 16559 7098
rect 16583 7046 16597 7098
rect 16597 7046 16609 7098
rect 16609 7046 16639 7098
rect 16663 7046 16673 7098
rect 16673 7046 16719 7098
rect 16423 7044 16479 7046
rect 16503 7044 16559 7046
rect 16583 7044 16639 7046
rect 16663 7044 16719 7046
rect 16423 6010 16479 6012
rect 16503 6010 16559 6012
rect 16583 6010 16639 6012
rect 16663 6010 16719 6012
rect 16423 5958 16469 6010
rect 16469 5958 16479 6010
rect 16503 5958 16533 6010
rect 16533 5958 16545 6010
rect 16545 5958 16559 6010
rect 16583 5958 16597 6010
rect 16597 5958 16609 6010
rect 16609 5958 16639 6010
rect 16663 5958 16673 6010
rect 16673 5958 16719 6010
rect 16423 5956 16479 5958
rect 16503 5956 16559 5958
rect 16583 5956 16639 5958
rect 16663 5956 16719 5958
rect 16302 5616 16358 5672
rect 16026 5228 16082 5264
rect 16026 5208 16028 5228
rect 16028 5208 16080 5228
rect 16080 5208 16082 5228
rect 16423 4922 16479 4924
rect 16503 4922 16559 4924
rect 16583 4922 16639 4924
rect 16663 4922 16719 4924
rect 16423 4870 16469 4922
rect 16469 4870 16479 4922
rect 16503 4870 16533 4922
rect 16533 4870 16545 4922
rect 16545 4870 16559 4922
rect 16583 4870 16597 4922
rect 16597 4870 16609 4922
rect 16609 4870 16639 4922
rect 16663 4870 16673 4922
rect 16673 4870 16719 4922
rect 16423 4868 16479 4870
rect 16503 4868 16559 4870
rect 16583 4868 16639 4870
rect 16663 4868 16719 4870
rect 16394 4700 16396 4720
rect 16396 4700 16448 4720
rect 16448 4700 16450 4720
rect 16394 4664 16450 4700
rect 16423 3834 16479 3836
rect 16503 3834 16559 3836
rect 16583 3834 16639 3836
rect 16663 3834 16719 3836
rect 16423 3782 16469 3834
rect 16469 3782 16479 3834
rect 16503 3782 16533 3834
rect 16533 3782 16545 3834
rect 16545 3782 16559 3834
rect 16583 3782 16597 3834
rect 16597 3782 16609 3834
rect 16609 3782 16639 3834
rect 16663 3782 16673 3834
rect 16673 3782 16719 3834
rect 16423 3780 16479 3782
rect 16503 3780 16559 3782
rect 16583 3780 16639 3782
rect 16663 3780 16719 3782
rect 17038 9632 17094 9688
rect 17774 9832 17830 9888
rect 17682 9632 17738 9688
rect 17083 8730 17139 8732
rect 17163 8730 17219 8732
rect 17243 8730 17299 8732
rect 17323 8730 17379 8732
rect 17083 8678 17129 8730
rect 17129 8678 17139 8730
rect 17163 8678 17193 8730
rect 17193 8678 17205 8730
rect 17205 8678 17219 8730
rect 17243 8678 17257 8730
rect 17257 8678 17269 8730
rect 17269 8678 17299 8730
rect 17323 8678 17333 8730
rect 17333 8678 17379 8730
rect 17083 8676 17139 8678
rect 17163 8676 17219 8678
rect 17243 8676 17299 8678
rect 17323 8676 17379 8678
rect 17083 7642 17139 7644
rect 17163 7642 17219 7644
rect 17243 7642 17299 7644
rect 17323 7642 17379 7644
rect 17083 7590 17129 7642
rect 17129 7590 17139 7642
rect 17163 7590 17193 7642
rect 17193 7590 17205 7642
rect 17205 7590 17219 7642
rect 17243 7590 17257 7642
rect 17257 7590 17269 7642
rect 17269 7590 17299 7642
rect 17323 7590 17333 7642
rect 17333 7590 17379 7642
rect 17083 7588 17139 7590
rect 17163 7588 17219 7590
rect 17243 7588 17299 7590
rect 17323 7588 17379 7590
rect 17083 6554 17139 6556
rect 17163 6554 17219 6556
rect 17243 6554 17299 6556
rect 17323 6554 17379 6556
rect 17083 6502 17129 6554
rect 17129 6502 17139 6554
rect 17163 6502 17193 6554
rect 17193 6502 17205 6554
rect 17205 6502 17219 6554
rect 17243 6502 17257 6554
rect 17257 6502 17269 6554
rect 17269 6502 17299 6554
rect 17323 6502 17333 6554
rect 17333 6502 17379 6554
rect 17083 6500 17139 6502
rect 17163 6500 17219 6502
rect 17243 6500 17299 6502
rect 17323 6500 17379 6502
rect 17130 5652 17132 5672
rect 17132 5652 17184 5672
rect 17184 5652 17186 5672
rect 17130 5616 17186 5652
rect 17083 5466 17139 5468
rect 17163 5466 17219 5468
rect 17243 5466 17299 5468
rect 17323 5466 17379 5468
rect 17083 5414 17129 5466
rect 17129 5414 17139 5466
rect 17163 5414 17193 5466
rect 17193 5414 17205 5466
rect 17205 5414 17219 5466
rect 17243 5414 17257 5466
rect 17257 5414 17269 5466
rect 17269 5414 17299 5466
rect 17323 5414 17333 5466
rect 17333 5414 17379 5466
rect 17083 5412 17139 5414
rect 17163 5412 17219 5414
rect 17243 5412 17299 5414
rect 17323 5412 17379 5414
rect 16423 2746 16479 2748
rect 16503 2746 16559 2748
rect 16583 2746 16639 2748
rect 16663 2746 16719 2748
rect 16423 2694 16469 2746
rect 16469 2694 16479 2746
rect 16503 2694 16533 2746
rect 16533 2694 16545 2746
rect 16545 2694 16559 2746
rect 16583 2694 16597 2746
rect 16597 2694 16609 2746
rect 16609 2694 16639 2746
rect 16663 2694 16673 2746
rect 16673 2694 16719 2746
rect 16423 2692 16479 2694
rect 16503 2692 16559 2694
rect 16583 2692 16639 2694
rect 16663 2692 16719 2694
rect 17083 4378 17139 4380
rect 17163 4378 17219 4380
rect 17243 4378 17299 4380
rect 17323 4378 17379 4380
rect 17083 4326 17129 4378
rect 17129 4326 17139 4378
rect 17163 4326 17193 4378
rect 17193 4326 17205 4378
rect 17205 4326 17219 4378
rect 17243 4326 17257 4378
rect 17257 4326 17269 4378
rect 17269 4326 17299 4378
rect 17323 4326 17333 4378
rect 17333 4326 17379 4378
rect 17083 4324 17139 4326
rect 17163 4324 17219 4326
rect 17243 4324 17299 4326
rect 17323 4324 17379 4326
rect 17083 3290 17139 3292
rect 17163 3290 17219 3292
rect 17243 3290 17299 3292
rect 17323 3290 17379 3292
rect 17083 3238 17129 3290
rect 17129 3238 17139 3290
rect 17163 3238 17193 3290
rect 17193 3238 17205 3290
rect 17205 3238 17219 3290
rect 17243 3238 17257 3290
rect 17257 3238 17269 3290
rect 17269 3238 17299 3290
rect 17323 3238 17333 3290
rect 17333 3238 17379 3290
rect 17083 3236 17139 3238
rect 17163 3236 17219 3238
rect 17243 3236 17299 3238
rect 17323 3236 17379 3238
rect 17682 7248 17738 7304
rect 17774 6568 17830 6624
rect 17958 6296 18014 6352
rect 19614 10104 19670 10160
rect 21546 17992 21602 18048
rect 20534 13252 20590 13288
rect 20534 13232 20536 13252
rect 20536 13232 20588 13252
rect 20588 13232 20590 13252
rect 20718 10648 20774 10704
rect 21086 4528 21142 4584
rect 21086 3032 21142 3088
rect 25502 27920 25558 27976
rect 24858 26560 24914 26616
rect 22610 25594 22666 25596
rect 22690 25594 22746 25596
rect 22770 25594 22826 25596
rect 22850 25594 22906 25596
rect 22610 25542 22656 25594
rect 22656 25542 22666 25594
rect 22690 25542 22720 25594
rect 22720 25542 22732 25594
rect 22732 25542 22746 25594
rect 22770 25542 22784 25594
rect 22784 25542 22796 25594
rect 22796 25542 22826 25594
rect 22850 25542 22860 25594
rect 22860 25542 22906 25594
rect 22610 25540 22666 25542
rect 22690 25540 22746 25542
rect 22770 25540 22826 25542
rect 22850 25540 22906 25542
rect 22610 24506 22666 24508
rect 22690 24506 22746 24508
rect 22770 24506 22826 24508
rect 22850 24506 22906 24508
rect 22610 24454 22656 24506
rect 22656 24454 22666 24506
rect 22690 24454 22720 24506
rect 22720 24454 22732 24506
rect 22732 24454 22746 24506
rect 22770 24454 22784 24506
rect 22784 24454 22796 24506
rect 22796 24454 22826 24506
rect 22850 24454 22860 24506
rect 22860 24454 22906 24506
rect 22610 24452 22666 24454
rect 22690 24452 22746 24454
rect 22770 24452 22826 24454
rect 22850 24452 22906 24454
rect 22610 23418 22666 23420
rect 22690 23418 22746 23420
rect 22770 23418 22826 23420
rect 22850 23418 22906 23420
rect 22610 23366 22656 23418
rect 22656 23366 22666 23418
rect 22690 23366 22720 23418
rect 22720 23366 22732 23418
rect 22732 23366 22746 23418
rect 22770 23366 22784 23418
rect 22784 23366 22796 23418
rect 22796 23366 22826 23418
rect 22850 23366 22860 23418
rect 22860 23366 22906 23418
rect 22610 23364 22666 23366
rect 22690 23364 22746 23366
rect 22770 23364 22826 23366
rect 22850 23364 22906 23366
rect 22610 22330 22666 22332
rect 22690 22330 22746 22332
rect 22770 22330 22826 22332
rect 22850 22330 22906 22332
rect 22610 22278 22656 22330
rect 22656 22278 22666 22330
rect 22690 22278 22720 22330
rect 22720 22278 22732 22330
rect 22732 22278 22746 22330
rect 22770 22278 22784 22330
rect 22784 22278 22796 22330
rect 22796 22278 22826 22330
rect 22850 22278 22860 22330
rect 22860 22278 22906 22330
rect 22610 22276 22666 22278
rect 22690 22276 22746 22278
rect 22770 22276 22826 22278
rect 22850 22276 22906 22278
rect 22610 21242 22666 21244
rect 22690 21242 22746 21244
rect 22770 21242 22826 21244
rect 22850 21242 22906 21244
rect 22610 21190 22656 21242
rect 22656 21190 22666 21242
rect 22690 21190 22720 21242
rect 22720 21190 22732 21242
rect 22732 21190 22746 21242
rect 22770 21190 22784 21242
rect 22784 21190 22796 21242
rect 22796 21190 22826 21242
rect 22850 21190 22860 21242
rect 22860 21190 22906 21242
rect 22610 21188 22666 21190
rect 22690 21188 22746 21190
rect 22770 21188 22826 21190
rect 22850 21188 22906 21190
rect 22610 20154 22666 20156
rect 22690 20154 22746 20156
rect 22770 20154 22826 20156
rect 22850 20154 22906 20156
rect 22610 20102 22656 20154
rect 22656 20102 22666 20154
rect 22690 20102 22720 20154
rect 22720 20102 22732 20154
rect 22732 20102 22746 20154
rect 22770 20102 22784 20154
rect 22784 20102 22796 20154
rect 22796 20102 22826 20154
rect 22850 20102 22860 20154
rect 22860 20102 22906 20154
rect 22610 20100 22666 20102
rect 22690 20100 22746 20102
rect 22770 20100 22826 20102
rect 22850 20100 22906 20102
rect 22610 19066 22666 19068
rect 22690 19066 22746 19068
rect 22770 19066 22826 19068
rect 22850 19066 22906 19068
rect 22610 19014 22656 19066
rect 22656 19014 22666 19066
rect 22690 19014 22720 19066
rect 22720 19014 22732 19066
rect 22732 19014 22746 19066
rect 22770 19014 22784 19066
rect 22784 19014 22796 19066
rect 22796 19014 22826 19066
rect 22850 19014 22860 19066
rect 22860 19014 22906 19066
rect 22610 19012 22666 19014
rect 22690 19012 22746 19014
rect 22770 19012 22826 19014
rect 22850 19012 22906 19014
rect 22610 17978 22666 17980
rect 22690 17978 22746 17980
rect 22770 17978 22826 17980
rect 22850 17978 22906 17980
rect 22610 17926 22656 17978
rect 22656 17926 22666 17978
rect 22690 17926 22720 17978
rect 22720 17926 22732 17978
rect 22732 17926 22746 17978
rect 22770 17926 22784 17978
rect 22784 17926 22796 17978
rect 22796 17926 22826 17978
rect 22850 17926 22860 17978
rect 22860 17926 22906 17978
rect 22610 17924 22666 17926
rect 22690 17924 22746 17926
rect 22770 17924 22826 17926
rect 22850 17924 22906 17926
rect 22610 16890 22666 16892
rect 22690 16890 22746 16892
rect 22770 16890 22826 16892
rect 22850 16890 22906 16892
rect 22610 16838 22656 16890
rect 22656 16838 22666 16890
rect 22690 16838 22720 16890
rect 22720 16838 22732 16890
rect 22732 16838 22746 16890
rect 22770 16838 22784 16890
rect 22784 16838 22796 16890
rect 22796 16838 22826 16890
rect 22850 16838 22860 16890
rect 22860 16838 22906 16890
rect 22610 16836 22666 16838
rect 22690 16836 22746 16838
rect 22770 16836 22826 16838
rect 22850 16836 22906 16838
rect 22374 15952 22430 16008
rect 22610 15802 22666 15804
rect 22690 15802 22746 15804
rect 22770 15802 22826 15804
rect 22850 15802 22906 15804
rect 22610 15750 22656 15802
rect 22656 15750 22666 15802
rect 22690 15750 22720 15802
rect 22720 15750 22732 15802
rect 22732 15750 22746 15802
rect 22770 15750 22784 15802
rect 22784 15750 22796 15802
rect 22796 15750 22826 15802
rect 22850 15750 22860 15802
rect 22860 15750 22906 15802
rect 22610 15748 22666 15750
rect 22690 15748 22746 15750
rect 22770 15748 22826 15750
rect 22850 15748 22906 15750
rect 23270 26138 23326 26140
rect 23350 26138 23406 26140
rect 23430 26138 23486 26140
rect 23510 26138 23566 26140
rect 23270 26086 23316 26138
rect 23316 26086 23326 26138
rect 23350 26086 23380 26138
rect 23380 26086 23392 26138
rect 23392 26086 23406 26138
rect 23430 26086 23444 26138
rect 23444 26086 23456 26138
rect 23456 26086 23486 26138
rect 23510 26086 23520 26138
rect 23520 26086 23566 26138
rect 23270 26084 23326 26086
rect 23350 26084 23406 26086
rect 23430 26084 23486 26086
rect 23510 26084 23566 26086
rect 23270 25050 23326 25052
rect 23350 25050 23406 25052
rect 23430 25050 23486 25052
rect 23510 25050 23566 25052
rect 23270 24998 23316 25050
rect 23316 24998 23326 25050
rect 23350 24998 23380 25050
rect 23380 24998 23392 25050
rect 23392 24998 23406 25050
rect 23430 24998 23444 25050
rect 23444 24998 23456 25050
rect 23456 24998 23486 25050
rect 23510 24998 23520 25050
rect 23520 24998 23566 25050
rect 23270 24996 23326 24998
rect 23350 24996 23406 24998
rect 23430 24996 23486 24998
rect 23510 24996 23566 24998
rect 23270 23962 23326 23964
rect 23350 23962 23406 23964
rect 23430 23962 23486 23964
rect 23510 23962 23566 23964
rect 23270 23910 23316 23962
rect 23316 23910 23326 23962
rect 23350 23910 23380 23962
rect 23380 23910 23392 23962
rect 23392 23910 23406 23962
rect 23430 23910 23444 23962
rect 23444 23910 23456 23962
rect 23456 23910 23486 23962
rect 23510 23910 23520 23962
rect 23520 23910 23566 23962
rect 23270 23908 23326 23910
rect 23350 23908 23406 23910
rect 23430 23908 23486 23910
rect 23510 23908 23566 23910
rect 23270 22874 23326 22876
rect 23350 22874 23406 22876
rect 23430 22874 23486 22876
rect 23510 22874 23566 22876
rect 23270 22822 23316 22874
rect 23316 22822 23326 22874
rect 23350 22822 23380 22874
rect 23380 22822 23392 22874
rect 23392 22822 23406 22874
rect 23430 22822 23444 22874
rect 23444 22822 23456 22874
rect 23456 22822 23486 22874
rect 23510 22822 23520 22874
rect 23520 22822 23566 22874
rect 23270 22820 23326 22822
rect 23350 22820 23406 22822
rect 23430 22820 23486 22822
rect 23510 22820 23566 22822
rect 25318 25900 25374 25936
rect 25318 25880 25320 25900
rect 25320 25880 25372 25900
rect 25372 25880 25374 25900
rect 23270 21786 23326 21788
rect 23350 21786 23406 21788
rect 23430 21786 23486 21788
rect 23510 21786 23566 21788
rect 23270 21734 23316 21786
rect 23316 21734 23326 21786
rect 23350 21734 23380 21786
rect 23380 21734 23392 21786
rect 23392 21734 23406 21786
rect 23430 21734 23444 21786
rect 23444 21734 23456 21786
rect 23456 21734 23486 21786
rect 23510 21734 23520 21786
rect 23520 21734 23566 21786
rect 23270 21732 23326 21734
rect 23350 21732 23406 21734
rect 23430 21732 23486 21734
rect 23510 21732 23566 21734
rect 23270 20698 23326 20700
rect 23350 20698 23406 20700
rect 23430 20698 23486 20700
rect 23510 20698 23566 20700
rect 23270 20646 23316 20698
rect 23316 20646 23326 20698
rect 23350 20646 23380 20698
rect 23380 20646 23392 20698
rect 23392 20646 23406 20698
rect 23430 20646 23444 20698
rect 23444 20646 23456 20698
rect 23456 20646 23486 20698
rect 23510 20646 23520 20698
rect 23520 20646 23566 20698
rect 23270 20644 23326 20646
rect 23350 20644 23406 20646
rect 23430 20644 23486 20646
rect 23510 20644 23566 20646
rect 23270 19610 23326 19612
rect 23350 19610 23406 19612
rect 23430 19610 23486 19612
rect 23510 19610 23566 19612
rect 23270 19558 23316 19610
rect 23316 19558 23326 19610
rect 23350 19558 23380 19610
rect 23380 19558 23392 19610
rect 23392 19558 23406 19610
rect 23430 19558 23444 19610
rect 23444 19558 23456 19610
rect 23456 19558 23486 19610
rect 23510 19558 23520 19610
rect 23520 19558 23566 19610
rect 23270 19556 23326 19558
rect 23350 19556 23406 19558
rect 23430 19556 23486 19558
rect 23510 19556 23566 19558
rect 23270 18522 23326 18524
rect 23350 18522 23406 18524
rect 23430 18522 23486 18524
rect 23510 18522 23566 18524
rect 23270 18470 23316 18522
rect 23316 18470 23326 18522
rect 23350 18470 23380 18522
rect 23380 18470 23392 18522
rect 23392 18470 23406 18522
rect 23430 18470 23444 18522
rect 23444 18470 23456 18522
rect 23456 18470 23486 18522
rect 23510 18470 23520 18522
rect 23520 18470 23566 18522
rect 23270 18468 23326 18470
rect 23350 18468 23406 18470
rect 23430 18468 23486 18470
rect 23510 18468 23566 18470
rect 23270 17434 23326 17436
rect 23350 17434 23406 17436
rect 23430 17434 23486 17436
rect 23510 17434 23566 17436
rect 23270 17382 23316 17434
rect 23316 17382 23326 17434
rect 23350 17382 23380 17434
rect 23380 17382 23392 17434
rect 23392 17382 23406 17434
rect 23430 17382 23444 17434
rect 23444 17382 23456 17434
rect 23456 17382 23486 17434
rect 23510 17382 23520 17434
rect 23520 17382 23566 17434
rect 23270 17380 23326 17382
rect 23350 17380 23406 17382
rect 23430 17380 23486 17382
rect 23510 17380 23566 17382
rect 23270 16346 23326 16348
rect 23350 16346 23406 16348
rect 23430 16346 23486 16348
rect 23510 16346 23566 16348
rect 23270 16294 23316 16346
rect 23316 16294 23326 16346
rect 23350 16294 23380 16346
rect 23380 16294 23392 16346
rect 23392 16294 23406 16346
rect 23430 16294 23444 16346
rect 23444 16294 23456 16346
rect 23456 16294 23486 16346
rect 23510 16294 23520 16346
rect 23520 16294 23566 16346
rect 23270 16292 23326 16294
rect 23350 16292 23406 16294
rect 23430 16292 23486 16294
rect 23510 16292 23566 16294
rect 23202 16108 23258 16144
rect 23202 16088 23204 16108
rect 23204 16088 23256 16108
rect 23256 16088 23258 16108
rect 23386 16088 23442 16144
rect 23846 19780 23902 19816
rect 23846 19760 23848 19780
rect 23848 19760 23900 19780
rect 23900 19760 23902 19780
rect 23270 15258 23326 15260
rect 23350 15258 23406 15260
rect 23430 15258 23486 15260
rect 23510 15258 23566 15260
rect 23270 15206 23316 15258
rect 23316 15206 23326 15258
rect 23350 15206 23380 15258
rect 23380 15206 23392 15258
rect 23392 15206 23406 15258
rect 23430 15206 23444 15258
rect 23444 15206 23456 15258
rect 23456 15206 23486 15258
rect 23510 15206 23520 15258
rect 23520 15206 23566 15258
rect 23270 15204 23326 15206
rect 23350 15204 23406 15206
rect 23430 15204 23486 15206
rect 23510 15204 23566 15206
rect 22190 14320 22246 14376
rect 22610 14714 22666 14716
rect 22690 14714 22746 14716
rect 22770 14714 22826 14716
rect 22850 14714 22906 14716
rect 22610 14662 22656 14714
rect 22656 14662 22666 14714
rect 22690 14662 22720 14714
rect 22720 14662 22732 14714
rect 22732 14662 22746 14714
rect 22770 14662 22784 14714
rect 22784 14662 22796 14714
rect 22796 14662 22826 14714
rect 22850 14662 22860 14714
rect 22860 14662 22906 14714
rect 22610 14660 22666 14662
rect 22690 14660 22746 14662
rect 22770 14660 22826 14662
rect 22850 14660 22906 14662
rect 22610 13626 22666 13628
rect 22690 13626 22746 13628
rect 22770 13626 22826 13628
rect 22850 13626 22906 13628
rect 22610 13574 22656 13626
rect 22656 13574 22666 13626
rect 22690 13574 22720 13626
rect 22720 13574 22732 13626
rect 22732 13574 22746 13626
rect 22770 13574 22784 13626
rect 22784 13574 22796 13626
rect 22796 13574 22826 13626
rect 22850 13574 22860 13626
rect 22860 13574 22906 13626
rect 22610 13572 22666 13574
rect 22690 13572 22746 13574
rect 22770 13572 22826 13574
rect 22850 13572 22906 13574
rect 22610 12538 22666 12540
rect 22690 12538 22746 12540
rect 22770 12538 22826 12540
rect 22850 12538 22906 12540
rect 22610 12486 22656 12538
rect 22656 12486 22666 12538
rect 22690 12486 22720 12538
rect 22720 12486 22732 12538
rect 22732 12486 22746 12538
rect 22770 12486 22784 12538
rect 22784 12486 22796 12538
rect 22796 12486 22826 12538
rect 22850 12486 22860 12538
rect 22860 12486 22906 12538
rect 22610 12484 22666 12486
rect 22690 12484 22746 12486
rect 22770 12484 22826 12486
rect 22850 12484 22906 12486
rect 22610 11450 22666 11452
rect 22690 11450 22746 11452
rect 22770 11450 22826 11452
rect 22850 11450 22906 11452
rect 22610 11398 22656 11450
rect 22656 11398 22666 11450
rect 22690 11398 22720 11450
rect 22720 11398 22732 11450
rect 22732 11398 22746 11450
rect 22770 11398 22784 11450
rect 22784 11398 22796 11450
rect 22796 11398 22826 11450
rect 22850 11398 22860 11450
rect 22860 11398 22906 11450
rect 22610 11396 22666 11398
rect 22690 11396 22746 11398
rect 22770 11396 22826 11398
rect 22850 11396 22906 11398
rect 23270 14170 23326 14172
rect 23350 14170 23406 14172
rect 23430 14170 23486 14172
rect 23510 14170 23566 14172
rect 23270 14118 23316 14170
rect 23316 14118 23326 14170
rect 23350 14118 23380 14170
rect 23380 14118 23392 14170
rect 23392 14118 23406 14170
rect 23430 14118 23444 14170
rect 23444 14118 23456 14170
rect 23456 14118 23486 14170
rect 23510 14118 23520 14170
rect 23520 14118 23566 14170
rect 23270 14116 23326 14118
rect 23350 14116 23406 14118
rect 23430 14116 23486 14118
rect 23510 14116 23566 14118
rect 23270 13082 23326 13084
rect 23350 13082 23406 13084
rect 23430 13082 23486 13084
rect 23510 13082 23566 13084
rect 23270 13030 23316 13082
rect 23316 13030 23326 13082
rect 23350 13030 23380 13082
rect 23380 13030 23392 13082
rect 23392 13030 23406 13082
rect 23430 13030 23444 13082
rect 23444 13030 23456 13082
rect 23456 13030 23486 13082
rect 23510 13030 23520 13082
rect 23520 13030 23566 13082
rect 23270 13028 23326 13030
rect 23350 13028 23406 13030
rect 23430 13028 23486 13030
rect 23510 13028 23566 13030
rect 22610 10362 22666 10364
rect 22690 10362 22746 10364
rect 22770 10362 22826 10364
rect 22850 10362 22906 10364
rect 22610 10310 22656 10362
rect 22656 10310 22666 10362
rect 22690 10310 22720 10362
rect 22720 10310 22732 10362
rect 22732 10310 22746 10362
rect 22770 10310 22784 10362
rect 22784 10310 22796 10362
rect 22796 10310 22826 10362
rect 22850 10310 22860 10362
rect 22860 10310 22906 10362
rect 22610 10308 22666 10310
rect 22690 10308 22746 10310
rect 22770 10308 22826 10310
rect 22850 10308 22906 10310
rect 23938 15408 23994 15464
rect 23270 11994 23326 11996
rect 23350 11994 23406 11996
rect 23430 11994 23486 11996
rect 23510 11994 23566 11996
rect 23270 11942 23316 11994
rect 23316 11942 23326 11994
rect 23350 11942 23380 11994
rect 23380 11942 23392 11994
rect 23392 11942 23406 11994
rect 23430 11942 23444 11994
rect 23444 11942 23456 11994
rect 23456 11942 23486 11994
rect 23510 11942 23520 11994
rect 23520 11942 23566 11994
rect 23270 11940 23326 11942
rect 23350 11940 23406 11942
rect 23430 11940 23486 11942
rect 23510 11940 23566 11942
rect 23270 10906 23326 10908
rect 23350 10906 23406 10908
rect 23430 10906 23486 10908
rect 23510 10906 23566 10908
rect 23270 10854 23316 10906
rect 23316 10854 23326 10906
rect 23350 10854 23380 10906
rect 23380 10854 23392 10906
rect 23392 10854 23406 10906
rect 23430 10854 23444 10906
rect 23444 10854 23456 10906
rect 23456 10854 23486 10906
rect 23510 10854 23520 10906
rect 23520 10854 23566 10906
rect 23270 10852 23326 10854
rect 23350 10852 23406 10854
rect 23430 10852 23486 10854
rect 23510 10852 23566 10854
rect 2778 720 2834 776
rect 19430 2352 19486 2408
rect 17083 2202 17139 2204
rect 17163 2202 17219 2204
rect 17243 2202 17299 2204
rect 17323 2202 17379 2204
rect 17083 2150 17129 2202
rect 17129 2150 17139 2202
rect 17163 2150 17193 2202
rect 17193 2150 17205 2202
rect 17205 2150 17219 2202
rect 17243 2150 17257 2202
rect 17257 2150 17269 2202
rect 17269 2150 17299 2202
rect 17323 2150 17333 2202
rect 17333 2150 17379 2202
rect 17083 2148 17139 2150
rect 17163 2148 17219 2150
rect 17243 2148 17299 2150
rect 17323 2148 17379 2150
rect 22610 9274 22666 9276
rect 22690 9274 22746 9276
rect 22770 9274 22826 9276
rect 22850 9274 22906 9276
rect 22610 9222 22656 9274
rect 22656 9222 22666 9274
rect 22690 9222 22720 9274
rect 22720 9222 22732 9274
rect 22732 9222 22746 9274
rect 22770 9222 22784 9274
rect 22784 9222 22796 9274
rect 22796 9222 22826 9274
rect 22850 9222 22860 9274
rect 22860 9222 22906 9274
rect 22610 9220 22666 9222
rect 22690 9220 22746 9222
rect 22770 9220 22826 9222
rect 22850 9220 22906 9222
rect 22610 8186 22666 8188
rect 22690 8186 22746 8188
rect 22770 8186 22826 8188
rect 22850 8186 22906 8188
rect 22610 8134 22656 8186
rect 22656 8134 22666 8186
rect 22690 8134 22720 8186
rect 22720 8134 22732 8186
rect 22732 8134 22746 8186
rect 22770 8134 22784 8186
rect 22784 8134 22796 8186
rect 22796 8134 22826 8186
rect 22850 8134 22860 8186
rect 22860 8134 22906 8186
rect 22610 8132 22666 8134
rect 22690 8132 22746 8134
rect 22770 8132 22826 8134
rect 22850 8132 22906 8134
rect 22610 7098 22666 7100
rect 22690 7098 22746 7100
rect 22770 7098 22826 7100
rect 22850 7098 22906 7100
rect 22610 7046 22656 7098
rect 22656 7046 22666 7098
rect 22690 7046 22720 7098
rect 22720 7046 22732 7098
rect 22732 7046 22746 7098
rect 22770 7046 22784 7098
rect 22784 7046 22796 7098
rect 22796 7046 22826 7098
rect 22850 7046 22860 7098
rect 22860 7046 22906 7098
rect 22610 7044 22666 7046
rect 22690 7044 22746 7046
rect 22770 7044 22826 7046
rect 22850 7044 22906 7046
rect 23270 9818 23326 9820
rect 23350 9818 23406 9820
rect 23430 9818 23486 9820
rect 23510 9818 23566 9820
rect 23270 9766 23316 9818
rect 23316 9766 23326 9818
rect 23350 9766 23380 9818
rect 23380 9766 23392 9818
rect 23392 9766 23406 9818
rect 23430 9766 23444 9818
rect 23444 9766 23456 9818
rect 23456 9766 23486 9818
rect 23510 9766 23520 9818
rect 23520 9766 23566 9818
rect 23270 9764 23326 9766
rect 23350 9764 23406 9766
rect 23430 9764 23486 9766
rect 23510 9764 23566 9766
rect 23270 8730 23326 8732
rect 23350 8730 23406 8732
rect 23430 8730 23486 8732
rect 23510 8730 23566 8732
rect 23270 8678 23316 8730
rect 23316 8678 23326 8730
rect 23350 8678 23380 8730
rect 23380 8678 23392 8730
rect 23392 8678 23406 8730
rect 23430 8678 23444 8730
rect 23444 8678 23456 8730
rect 23456 8678 23486 8730
rect 23510 8678 23520 8730
rect 23520 8678 23566 8730
rect 23270 8676 23326 8678
rect 23350 8676 23406 8678
rect 23430 8676 23486 8678
rect 23510 8676 23566 8678
rect 23270 7642 23326 7644
rect 23350 7642 23406 7644
rect 23430 7642 23486 7644
rect 23510 7642 23566 7644
rect 23270 7590 23316 7642
rect 23316 7590 23326 7642
rect 23350 7590 23380 7642
rect 23380 7590 23392 7642
rect 23392 7590 23406 7642
rect 23430 7590 23444 7642
rect 23444 7590 23456 7642
rect 23456 7590 23486 7642
rect 23510 7590 23520 7642
rect 23520 7590 23566 7642
rect 23270 7588 23326 7590
rect 23350 7588 23406 7590
rect 23430 7588 23486 7590
rect 23510 7588 23566 7590
rect 23270 6554 23326 6556
rect 23350 6554 23406 6556
rect 23430 6554 23486 6556
rect 23510 6554 23566 6556
rect 23270 6502 23316 6554
rect 23316 6502 23326 6554
rect 23350 6502 23380 6554
rect 23380 6502 23392 6554
rect 23392 6502 23406 6554
rect 23430 6502 23444 6554
rect 23444 6502 23456 6554
rect 23456 6502 23486 6554
rect 23510 6502 23520 6554
rect 23520 6502 23566 6554
rect 23270 6500 23326 6502
rect 23350 6500 23406 6502
rect 23430 6500 23486 6502
rect 23510 6500 23566 6502
rect 24858 25200 24914 25256
rect 25410 23840 25466 23896
rect 25410 19080 25466 19136
rect 25226 18808 25282 18864
rect 25042 16088 25098 16144
rect 25410 15700 25466 15736
rect 25410 15680 25412 15700
rect 25412 15680 25464 15700
rect 25464 15680 25466 15700
rect 25410 12960 25466 13016
rect 25410 10240 25466 10296
rect 25778 23160 25834 23216
rect 25686 17076 25688 17096
rect 25688 17076 25740 17096
rect 25740 17076 25742 17096
rect 25686 17040 25742 17076
rect 25686 13640 25742 13696
rect 24950 9968 25006 10024
rect 22610 6010 22666 6012
rect 22690 6010 22746 6012
rect 22770 6010 22826 6012
rect 22850 6010 22906 6012
rect 22610 5958 22656 6010
rect 22656 5958 22666 6010
rect 22690 5958 22720 6010
rect 22720 5958 22732 6010
rect 22732 5958 22746 6010
rect 22770 5958 22784 6010
rect 22784 5958 22796 6010
rect 22796 5958 22826 6010
rect 22850 5958 22860 6010
rect 22860 5958 22906 6010
rect 22610 5956 22666 5958
rect 22690 5956 22746 5958
rect 22770 5956 22826 5958
rect 22850 5956 22906 5958
rect 22610 4922 22666 4924
rect 22690 4922 22746 4924
rect 22770 4922 22826 4924
rect 22850 4922 22906 4924
rect 22610 4870 22656 4922
rect 22656 4870 22666 4922
rect 22690 4870 22720 4922
rect 22720 4870 22732 4922
rect 22732 4870 22746 4922
rect 22770 4870 22784 4922
rect 22784 4870 22796 4922
rect 22796 4870 22826 4922
rect 22850 4870 22860 4922
rect 22860 4870 22906 4922
rect 22610 4868 22666 4870
rect 22690 4868 22746 4870
rect 22770 4868 22826 4870
rect 22850 4868 22906 4870
rect 22610 3834 22666 3836
rect 22690 3834 22746 3836
rect 22770 3834 22826 3836
rect 22850 3834 22906 3836
rect 22610 3782 22656 3834
rect 22656 3782 22666 3834
rect 22690 3782 22720 3834
rect 22720 3782 22732 3834
rect 22732 3782 22746 3834
rect 22770 3782 22784 3834
rect 22784 3782 22796 3834
rect 22796 3782 22826 3834
rect 22850 3782 22860 3834
rect 22860 3782 22906 3834
rect 22610 3780 22666 3782
rect 22690 3780 22746 3782
rect 22770 3780 22826 3782
rect 22850 3780 22906 3782
rect 23270 5466 23326 5468
rect 23350 5466 23406 5468
rect 23430 5466 23486 5468
rect 23510 5466 23566 5468
rect 23270 5414 23316 5466
rect 23316 5414 23326 5466
rect 23350 5414 23380 5466
rect 23380 5414 23392 5466
rect 23392 5414 23406 5466
rect 23430 5414 23444 5466
rect 23444 5414 23456 5466
rect 23456 5414 23486 5466
rect 23510 5414 23520 5466
rect 23520 5414 23566 5466
rect 23270 5412 23326 5414
rect 23350 5412 23406 5414
rect 23430 5412 23486 5414
rect 23510 5412 23566 5414
rect 23270 4378 23326 4380
rect 23350 4378 23406 4380
rect 23430 4378 23486 4380
rect 23510 4378 23566 4380
rect 23270 4326 23316 4378
rect 23316 4326 23326 4378
rect 23350 4326 23380 4378
rect 23380 4326 23392 4378
rect 23392 4326 23406 4378
rect 23430 4326 23444 4378
rect 23444 4326 23456 4378
rect 23456 4326 23486 4378
rect 23510 4326 23520 4378
rect 23520 4326 23566 4378
rect 23270 4324 23326 4326
rect 23350 4324 23406 4326
rect 23430 4324 23486 4326
rect 23510 4324 23566 4326
rect 25962 22516 25964 22536
rect 25964 22516 26016 22536
rect 26016 22516 26018 22536
rect 25962 22480 26018 22516
rect 25962 21800 26018 21856
rect 25962 20440 26018 20496
rect 25962 19760 26018 19816
rect 25962 18400 26018 18456
rect 25962 16360 26018 16416
rect 25962 14320 26018 14376
rect 26330 12688 26386 12744
rect 26054 12280 26110 12336
rect 25962 10920 26018 10976
rect 25962 9560 26018 9616
rect 25962 8200 26018 8256
rect 25686 7520 25742 7576
rect 25962 6840 26018 6896
rect 25410 6180 25466 6216
rect 25410 6160 25412 6180
rect 25412 6160 25464 6180
rect 25464 6160 25466 6180
rect 25410 4800 25466 4856
rect 25410 4120 25466 4176
rect 23270 3290 23326 3292
rect 23350 3290 23406 3292
rect 23430 3290 23486 3292
rect 23510 3290 23566 3292
rect 23270 3238 23316 3290
rect 23316 3238 23326 3290
rect 23350 3238 23380 3290
rect 23380 3238 23392 3290
rect 23392 3238 23406 3290
rect 23430 3238 23444 3290
rect 23444 3238 23456 3290
rect 23456 3238 23486 3290
rect 23510 3238 23520 3290
rect 23520 3238 23566 3290
rect 23270 3236 23326 3238
rect 23350 3236 23406 3238
rect 23430 3236 23486 3238
rect 23510 3236 23566 3238
rect 22610 2746 22666 2748
rect 22690 2746 22746 2748
rect 22770 2746 22826 2748
rect 22850 2746 22906 2748
rect 22610 2694 22656 2746
rect 22656 2694 22666 2746
rect 22690 2694 22720 2746
rect 22720 2694 22732 2746
rect 22732 2694 22746 2746
rect 22770 2694 22784 2746
rect 22784 2694 22796 2746
rect 22796 2694 22826 2746
rect 22850 2694 22860 2746
rect 22860 2694 22906 2746
rect 22610 2692 22666 2694
rect 22690 2692 22746 2694
rect 22770 2692 22826 2694
rect 22850 2692 22906 2694
rect 23270 2202 23326 2204
rect 23350 2202 23406 2204
rect 23430 2202 23486 2204
rect 23510 2202 23566 2204
rect 23270 2150 23316 2202
rect 23316 2150 23326 2202
rect 23350 2150 23380 2202
rect 23380 2150 23392 2202
rect 23392 2150 23406 2202
rect 23430 2150 23444 2202
rect 23444 2150 23456 2202
rect 23456 2150 23486 2202
rect 23510 2150 23520 2202
rect 23520 2150 23566 2202
rect 23270 2148 23326 2150
rect 23350 2148 23406 2150
rect 23430 2148 23486 2150
rect 23510 2148 23566 2150
rect 25962 3476 25964 3496
rect 25964 3476 26016 3496
rect 26016 3476 26018 3496
rect 25962 3440 26018 3476
rect 25134 2796 25136 2816
rect 25136 2796 25188 2816
rect 25188 2796 25190 2816
rect 25134 2760 25190 2796
rect 24674 1400 24730 1456
rect 25042 856 25098 912
rect 25870 40 25926 96
<< metal3 >>
rect 0 28658 800 28688
rect 1577 28658 1643 28661
rect 0 28656 1643 28658
rect 0 28600 1582 28656
rect 1638 28600 1643 28656
rect 0 28598 1643 28600
rect 0 28568 800 28598
rect 1577 28595 1643 28598
rect 22921 28658 22987 28661
rect 26237 28658 27037 28688
rect 22921 28656 27037 28658
rect 22921 28600 22926 28656
rect 22982 28600 27037 28656
rect 22921 28598 27037 28600
rect 22921 28595 22987 28598
rect 26237 28568 27037 28598
rect 25497 27978 25563 27981
rect 26237 27978 27037 28008
rect 25497 27976 27037 27978
rect 25497 27920 25502 27976
rect 25558 27920 27037 27976
rect 25497 27918 27037 27920
rect 25497 27915 25563 27918
rect 26237 27888 27037 27918
rect 0 27298 800 27328
rect 0 27208 858 27298
rect 798 27026 858 27208
rect 1393 27026 1459 27029
rect 798 27024 1459 27026
rect 798 26968 1398 27024
rect 1454 26968 1459 27024
rect 798 26966 1459 26968
rect 1393 26963 1459 26966
rect 4039 26688 4355 26689
rect 0 26618 800 26648
rect 4039 26624 4045 26688
rect 4109 26624 4125 26688
rect 4189 26624 4205 26688
rect 4269 26624 4285 26688
rect 4349 26624 4355 26688
rect 4039 26623 4355 26624
rect 10226 26688 10542 26689
rect 10226 26624 10232 26688
rect 10296 26624 10312 26688
rect 10376 26624 10392 26688
rect 10456 26624 10472 26688
rect 10536 26624 10542 26688
rect 10226 26623 10542 26624
rect 16413 26688 16729 26689
rect 16413 26624 16419 26688
rect 16483 26624 16499 26688
rect 16563 26624 16579 26688
rect 16643 26624 16659 26688
rect 16723 26624 16729 26688
rect 16413 26623 16729 26624
rect 22600 26688 22916 26689
rect 22600 26624 22606 26688
rect 22670 26624 22686 26688
rect 22750 26624 22766 26688
rect 22830 26624 22846 26688
rect 22910 26624 22916 26688
rect 22600 26623 22916 26624
rect 2865 26618 2931 26621
rect 0 26616 2931 26618
rect 0 26560 2870 26616
rect 2926 26560 2931 26616
rect 0 26558 2931 26560
rect 0 26528 800 26558
rect 2865 26555 2931 26558
rect 24853 26618 24919 26621
rect 26237 26618 27037 26648
rect 24853 26616 27037 26618
rect 24853 26560 24858 26616
rect 24914 26560 27037 26616
rect 24853 26558 27037 26560
rect 24853 26555 24919 26558
rect 26237 26528 27037 26558
rect 4699 26144 5015 26145
rect 4699 26080 4705 26144
rect 4769 26080 4785 26144
rect 4849 26080 4865 26144
rect 4929 26080 4945 26144
rect 5009 26080 5015 26144
rect 4699 26079 5015 26080
rect 10886 26144 11202 26145
rect 10886 26080 10892 26144
rect 10956 26080 10972 26144
rect 11036 26080 11052 26144
rect 11116 26080 11132 26144
rect 11196 26080 11202 26144
rect 10886 26079 11202 26080
rect 17073 26144 17389 26145
rect 17073 26080 17079 26144
rect 17143 26080 17159 26144
rect 17223 26080 17239 26144
rect 17303 26080 17319 26144
rect 17383 26080 17389 26144
rect 17073 26079 17389 26080
rect 23260 26144 23576 26145
rect 23260 26080 23266 26144
rect 23330 26080 23346 26144
rect 23410 26080 23426 26144
rect 23490 26080 23506 26144
rect 23570 26080 23576 26144
rect 23260 26079 23576 26080
rect 0 25938 800 25968
rect 1025 25938 1091 25941
rect 0 25936 1091 25938
rect 0 25880 1030 25936
rect 1086 25880 1091 25936
rect 0 25878 1091 25880
rect 0 25848 800 25878
rect 1025 25875 1091 25878
rect 25313 25938 25379 25941
rect 26237 25938 27037 25968
rect 25313 25936 27037 25938
rect 25313 25880 25318 25936
rect 25374 25880 27037 25936
rect 25313 25878 27037 25880
rect 25313 25875 25379 25878
rect 26237 25848 27037 25878
rect 8569 25802 8635 25805
rect 15837 25802 15903 25805
rect 8569 25800 15903 25802
rect 8569 25744 8574 25800
rect 8630 25744 15842 25800
rect 15898 25744 15903 25800
rect 8569 25742 15903 25744
rect 8569 25739 8635 25742
rect 15837 25739 15903 25742
rect 4039 25600 4355 25601
rect 4039 25536 4045 25600
rect 4109 25536 4125 25600
rect 4189 25536 4205 25600
rect 4269 25536 4285 25600
rect 4349 25536 4355 25600
rect 4039 25535 4355 25536
rect 10226 25600 10542 25601
rect 10226 25536 10232 25600
rect 10296 25536 10312 25600
rect 10376 25536 10392 25600
rect 10456 25536 10472 25600
rect 10536 25536 10542 25600
rect 10226 25535 10542 25536
rect 16413 25600 16729 25601
rect 16413 25536 16419 25600
rect 16483 25536 16499 25600
rect 16563 25536 16579 25600
rect 16643 25536 16659 25600
rect 16723 25536 16729 25600
rect 16413 25535 16729 25536
rect 22600 25600 22916 25601
rect 22600 25536 22606 25600
rect 22670 25536 22686 25600
rect 22750 25536 22766 25600
rect 22830 25536 22846 25600
rect 22910 25536 22916 25600
rect 22600 25535 22916 25536
rect 10409 25394 10475 25397
rect 18505 25394 18571 25397
rect 10409 25392 18571 25394
rect 10409 25336 10414 25392
rect 10470 25336 18510 25392
rect 18566 25336 18571 25392
rect 10409 25334 18571 25336
rect 10409 25331 10475 25334
rect 18505 25331 18571 25334
rect 0 25258 800 25288
rect 1025 25258 1091 25261
rect 0 25256 1091 25258
rect 0 25200 1030 25256
rect 1086 25200 1091 25256
rect 0 25198 1091 25200
rect 0 25168 800 25198
rect 1025 25195 1091 25198
rect 24853 25258 24919 25261
rect 26237 25258 27037 25288
rect 24853 25256 27037 25258
rect 24853 25200 24858 25256
rect 24914 25200 27037 25256
rect 24853 25198 27037 25200
rect 24853 25195 24919 25198
rect 26237 25168 27037 25198
rect 4699 25056 5015 25057
rect 4699 24992 4705 25056
rect 4769 24992 4785 25056
rect 4849 24992 4865 25056
rect 4929 24992 4945 25056
rect 5009 24992 5015 25056
rect 4699 24991 5015 24992
rect 10886 25056 11202 25057
rect 10886 24992 10892 25056
rect 10956 24992 10972 25056
rect 11036 24992 11052 25056
rect 11116 24992 11132 25056
rect 11196 24992 11202 25056
rect 10886 24991 11202 24992
rect 17073 25056 17389 25057
rect 17073 24992 17079 25056
rect 17143 24992 17159 25056
rect 17223 24992 17239 25056
rect 17303 24992 17319 25056
rect 17383 24992 17389 25056
rect 17073 24991 17389 24992
rect 23260 25056 23576 25057
rect 23260 24992 23266 25056
rect 23330 24992 23346 25056
rect 23410 24992 23426 25056
rect 23490 24992 23506 25056
rect 23570 24992 23576 25056
rect 23260 24991 23576 24992
rect 6821 24850 6887 24853
rect 21081 24850 21147 24853
rect 6821 24848 21147 24850
rect 6821 24792 6826 24848
rect 6882 24792 21086 24848
rect 21142 24792 21147 24848
rect 6821 24790 21147 24792
rect 6821 24787 6887 24790
rect 21081 24787 21147 24790
rect 9673 24714 9739 24717
rect 9806 24714 9812 24716
rect 9673 24712 9812 24714
rect 9673 24656 9678 24712
rect 9734 24656 9812 24712
rect 9673 24654 9812 24656
rect 9673 24651 9739 24654
rect 9806 24652 9812 24654
rect 9876 24652 9882 24716
rect 4039 24512 4355 24513
rect 4039 24448 4045 24512
rect 4109 24448 4125 24512
rect 4189 24448 4205 24512
rect 4269 24448 4285 24512
rect 4349 24448 4355 24512
rect 4039 24447 4355 24448
rect 10226 24512 10542 24513
rect 10226 24448 10232 24512
rect 10296 24448 10312 24512
rect 10376 24448 10392 24512
rect 10456 24448 10472 24512
rect 10536 24448 10542 24512
rect 10226 24447 10542 24448
rect 16413 24512 16729 24513
rect 16413 24448 16419 24512
rect 16483 24448 16499 24512
rect 16563 24448 16579 24512
rect 16643 24448 16659 24512
rect 16723 24448 16729 24512
rect 16413 24447 16729 24448
rect 22600 24512 22916 24513
rect 22600 24448 22606 24512
rect 22670 24448 22686 24512
rect 22750 24448 22766 24512
rect 22830 24448 22846 24512
rect 22910 24448 22916 24512
rect 22600 24447 22916 24448
rect 12157 24306 12223 24309
rect 16389 24306 16455 24309
rect 12157 24304 16455 24306
rect 12157 24248 12162 24304
rect 12218 24248 16394 24304
rect 16450 24248 16455 24304
rect 12157 24246 16455 24248
rect 12157 24243 12223 24246
rect 16389 24243 16455 24246
rect 14365 24170 14431 24173
rect 17493 24170 17559 24173
rect 14365 24168 17559 24170
rect 14365 24112 14370 24168
rect 14426 24112 17498 24168
rect 17554 24112 17559 24168
rect 14365 24110 17559 24112
rect 14365 24107 14431 24110
rect 17493 24107 17559 24110
rect 4699 23968 5015 23969
rect 0 23898 800 23928
rect 4699 23904 4705 23968
rect 4769 23904 4785 23968
rect 4849 23904 4865 23968
rect 4929 23904 4945 23968
rect 5009 23904 5015 23968
rect 4699 23903 5015 23904
rect 10886 23968 11202 23969
rect 10886 23904 10892 23968
rect 10956 23904 10972 23968
rect 11036 23904 11052 23968
rect 11116 23904 11132 23968
rect 11196 23904 11202 23968
rect 10886 23903 11202 23904
rect 17073 23968 17389 23969
rect 17073 23904 17079 23968
rect 17143 23904 17159 23968
rect 17223 23904 17239 23968
rect 17303 23904 17319 23968
rect 17383 23904 17389 23968
rect 17073 23903 17389 23904
rect 23260 23968 23576 23969
rect 23260 23904 23266 23968
rect 23330 23904 23346 23968
rect 23410 23904 23426 23968
rect 23490 23904 23506 23968
rect 23570 23904 23576 23968
rect 23260 23903 23576 23904
rect 933 23898 999 23901
rect 0 23896 999 23898
rect 0 23840 938 23896
rect 994 23840 999 23896
rect 0 23838 999 23840
rect 0 23808 800 23838
rect 933 23835 999 23838
rect 9765 23898 9831 23901
rect 10501 23898 10567 23901
rect 9765 23896 10567 23898
rect 9765 23840 9770 23896
rect 9826 23840 10506 23896
rect 10562 23840 10567 23896
rect 9765 23838 10567 23840
rect 9765 23835 9831 23838
rect 10501 23835 10567 23838
rect 25405 23898 25471 23901
rect 26237 23898 27037 23928
rect 25405 23896 27037 23898
rect 25405 23840 25410 23896
rect 25466 23840 27037 23896
rect 25405 23838 27037 23840
rect 25405 23835 25471 23838
rect 26237 23808 27037 23838
rect 8753 23762 8819 23765
rect 10133 23762 10199 23765
rect 14549 23762 14615 23765
rect 8753 23760 14615 23762
rect 8753 23704 8758 23760
rect 8814 23704 10138 23760
rect 10194 23704 14554 23760
rect 14610 23704 14615 23760
rect 8753 23702 14615 23704
rect 8753 23699 8819 23702
rect 10133 23699 10199 23702
rect 14549 23699 14615 23702
rect 1577 23626 1643 23629
rect 21265 23626 21331 23629
rect 1577 23624 21331 23626
rect 1577 23568 1582 23624
rect 1638 23568 21270 23624
rect 21326 23568 21331 23624
rect 1577 23566 21331 23568
rect 1577 23563 1643 23566
rect 21265 23563 21331 23566
rect 1393 23488 1459 23493
rect 1393 23432 1398 23488
rect 1454 23432 1459 23488
rect 1393 23427 1459 23432
rect 0 23218 800 23248
rect 1396 23218 1456 23427
rect 4039 23424 4355 23425
rect 4039 23360 4045 23424
rect 4109 23360 4125 23424
rect 4189 23360 4205 23424
rect 4269 23360 4285 23424
rect 4349 23360 4355 23424
rect 4039 23359 4355 23360
rect 10226 23424 10542 23425
rect 10226 23360 10232 23424
rect 10296 23360 10312 23424
rect 10376 23360 10392 23424
rect 10456 23360 10472 23424
rect 10536 23360 10542 23424
rect 10226 23359 10542 23360
rect 16413 23424 16729 23425
rect 16413 23360 16419 23424
rect 16483 23360 16499 23424
rect 16563 23360 16579 23424
rect 16643 23360 16659 23424
rect 16723 23360 16729 23424
rect 16413 23359 16729 23360
rect 22600 23424 22916 23425
rect 22600 23360 22606 23424
rect 22670 23360 22686 23424
rect 22750 23360 22766 23424
rect 22830 23360 22846 23424
rect 22910 23360 22916 23424
rect 22600 23359 22916 23360
rect 0 23158 1456 23218
rect 25773 23218 25839 23221
rect 26237 23218 27037 23248
rect 25773 23216 27037 23218
rect 25773 23160 25778 23216
rect 25834 23160 27037 23216
rect 25773 23158 27037 23160
rect 0 23128 800 23158
rect 25773 23155 25839 23158
rect 26237 23128 27037 23158
rect 4699 22880 5015 22881
rect 4699 22816 4705 22880
rect 4769 22816 4785 22880
rect 4849 22816 4865 22880
rect 4929 22816 4945 22880
rect 5009 22816 5015 22880
rect 4699 22815 5015 22816
rect 10886 22880 11202 22881
rect 10886 22816 10892 22880
rect 10956 22816 10972 22880
rect 11036 22816 11052 22880
rect 11116 22816 11132 22880
rect 11196 22816 11202 22880
rect 10886 22815 11202 22816
rect 17073 22880 17389 22881
rect 17073 22816 17079 22880
rect 17143 22816 17159 22880
rect 17223 22816 17239 22880
rect 17303 22816 17319 22880
rect 17383 22816 17389 22880
rect 17073 22815 17389 22816
rect 23260 22880 23576 22881
rect 23260 22816 23266 22880
rect 23330 22816 23346 22880
rect 23410 22816 23426 22880
rect 23490 22816 23506 22880
rect 23570 22816 23576 22880
rect 23260 22815 23576 22816
rect 9765 22812 9831 22813
rect 9765 22810 9812 22812
rect 9720 22808 9812 22810
rect 9720 22752 9770 22808
rect 9720 22750 9812 22752
rect 9765 22748 9812 22750
rect 9876 22748 9882 22812
rect 9765 22747 9831 22748
rect 0 22538 800 22568
rect 933 22538 999 22541
rect 0 22536 999 22538
rect 0 22480 938 22536
rect 994 22480 999 22536
rect 0 22478 999 22480
rect 0 22448 800 22478
rect 933 22475 999 22478
rect 25957 22538 26023 22541
rect 26237 22538 27037 22568
rect 25957 22536 27037 22538
rect 25957 22480 25962 22536
rect 26018 22480 27037 22536
rect 25957 22478 27037 22480
rect 25957 22475 26023 22478
rect 26237 22448 27037 22478
rect 4039 22336 4355 22337
rect 4039 22272 4045 22336
rect 4109 22272 4125 22336
rect 4189 22272 4205 22336
rect 4269 22272 4285 22336
rect 4349 22272 4355 22336
rect 4039 22271 4355 22272
rect 10226 22336 10542 22337
rect 10226 22272 10232 22336
rect 10296 22272 10312 22336
rect 10376 22272 10392 22336
rect 10456 22272 10472 22336
rect 10536 22272 10542 22336
rect 10226 22271 10542 22272
rect 16413 22336 16729 22337
rect 16413 22272 16419 22336
rect 16483 22272 16499 22336
rect 16563 22272 16579 22336
rect 16643 22272 16659 22336
rect 16723 22272 16729 22336
rect 16413 22271 16729 22272
rect 22600 22336 22916 22337
rect 22600 22272 22606 22336
rect 22670 22272 22686 22336
rect 22750 22272 22766 22336
rect 22830 22272 22846 22336
rect 22910 22272 22916 22336
rect 22600 22271 22916 22272
rect 9949 22130 10015 22133
rect 10225 22130 10291 22133
rect 9949 22128 10291 22130
rect 9949 22072 9954 22128
rect 10010 22072 10230 22128
rect 10286 22072 10291 22128
rect 9949 22070 10291 22072
rect 9949 22067 10015 22070
rect 10225 22067 10291 22070
rect 17585 22130 17651 22133
rect 17585 22128 17786 22130
rect 17585 22072 17590 22128
rect 17646 22072 17786 22128
rect 17585 22070 17786 22072
rect 17585 22067 17651 22070
rect 10777 21994 10843 21997
rect 2730 21992 10843 21994
rect 2730 21936 10782 21992
rect 10838 21936 10843 21992
rect 2730 21934 10843 21936
rect 17726 21994 17786 22070
rect 17861 21994 17927 21997
rect 17726 21992 17927 21994
rect 17726 21936 17866 21992
rect 17922 21936 17927 21992
rect 17726 21934 17927 21936
rect 2405 21450 2471 21453
rect 2730 21450 2790 21934
rect 10777 21931 10843 21934
rect 17861 21931 17927 21934
rect 25957 21858 26023 21861
rect 26237 21858 27037 21888
rect 25957 21856 27037 21858
rect 25957 21800 25962 21856
rect 26018 21800 27037 21856
rect 25957 21798 27037 21800
rect 25957 21795 26023 21798
rect 4699 21792 5015 21793
rect 4699 21728 4705 21792
rect 4769 21728 4785 21792
rect 4849 21728 4865 21792
rect 4929 21728 4945 21792
rect 5009 21728 5015 21792
rect 4699 21727 5015 21728
rect 10886 21792 11202 21793
rect 10886 21728 10892 21792
rect 10956 21728 10972 21792
rect 11036 21728 11052 21792
rect 11116 21728 11132 21792
rect 11196 21728 11202 21792
rect 10886 21727 11202 21728
rect 17073 21792 17389 21793
rect 17073 21728 17079 21792
rect 17143 21728 17159 21792
rect 17223 21728 17239 21792
rect 17303 21728 17319 21792
rect 17383 21728 17389 21792
rect 17073 21727 17389 21728
rect 23260 21792 23576 21793
rect 23260 21728 23266 21792
rect 23330 21728 23346 21792
rect 23410 21728 23426 21792
rect 23490 21728 23506 21792
rect 23570 21728 23576 21792
rect 26237 21768 27037 21798
rect 23260 21727 23576 21728
rect 10041 21586 10107 21589
rect 15193 21586 15259 21589
rect 10041 21584 15259 21586
rect 10041 21528 10046 21584
rect 10102 21528 15198 21584
rect 15254 21528 15259 21584
rect 10041 21526 15259 21528
rect 10041 21523 10107 21526
rect 15193 21523 15259 21526
rect 2405 21448 2790 21450
rect 2405 21392 2410 21448
rect 2466 21392 2790 21448
rect 2405 21390 2790 21392
rect 2405 21387 2471 21390
rect 4039 21248 4355 21249
rect 0 21178 800 21208
rect 4039 21184 4045 21248
rect 4109 21184 4125 21248
rect 4189 21184 4205 21248
rect 4269 21184 4285 21248
rect 4349 21184 4355 21248
rect 4039 21183 4355 21184
rect 10226 21248 10542 21249
rect 10226 21184 10232 21248
rect 10296 21184 10312 21248
rect 10376 21184 10392 21248
rect 10456 21184 10472 21248
rect 10536 21184 10542 21248
rect 10226 21183 10542 21184
rect 16413 21248 16729 21249
rect 16413 21184 16419 21248
rect 16483 21184 16499 21248
rect 16563 21184 16579 21248
rect 16643 21184 16659 21248
rect 16723 21184 16729 21248
rect 16413 21183 16729 21184
rect 22600 21248 22916 21249
rect 22600 21184 22606 21248
rect 22670 21184 22686 21248
rect 22750 21184 22766 21248
rect 22830 21184 22846 21248
rect 22910 21184 22916 21248
rect 22600 21183 22916 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 7833 20772 7899 20773
rect 7782 20708 7788 20772
rect 7852 20770 7899 20772
rect 7852 20768 7944 20770
rect 7894 20712 7944 20768
rect 7852 20710 7944 20712
rect 7852 20708 7899 20710
rect 7833 20707 7899 20708
rect 4699 20704 5015 20705
rect 4699 20640 4705 20704
rect 4769 20640 4785 20704
rect 4849 20640 4865 20704
rect 4929 20640 4945 20704
rect 5009 20640 5015 20704
rect 4699 20639 5015 20640
rect 10886 20704 11202 20705
rect 10886 20640 10892 20704
rect 10956 20640 10972 20704
rect 11036 20640 11052 20704
rect 11116 20640 11132 20704
rect 11196 20640 11202 20704
rect 10886 20639 11202 20640
rect 17073 20704 17389 20705
rect 17073 20640 17079 20704
rect 17143 20640 17159 20704
rect 17223 20640 17239 20704
rect 17303 20640 17319 20704
rect 17383 20640 17389 20704
rect 17073 20639 17389 20640
rect 23260 20704 23576 20705
rect 23260 20640 23266 20704
rect 23330 20640 23346 20704
rect 23410 20640 23426 20704
rect 23490 20640 23506 20704
rect 23570 20640 23576 20704
rect 23260 20639 23576 20640
rect 1393 20632 1459 20637
rect 1393 20576 1398 20632
rect 1454 20576 1459 20632
rect 1393 20571 1459 20576
rect 0 20498 800 20528
rect 1396 20498 1456 20571
rect 0 20438 1456 20498
rect 2681 20498 2747 20501
rect 25957 20498 26023 20501
rect 26237 20498 27037 20528
rect 2681 20496 2790 20498
rect 2681 20440 2686 20496
rect 2742 20440 2790 20496
rect 0 20408 800 20438
rect 2681 20435 2790 20440
rect 25957 20496 27037 20498
rect 25957 20440 25962 20496
rect 26018 20440 27037 20496
rect 25957 20438 27037 20440
rect 25957 20435 26023 20438
rect 0 19818 800 19848
rect 2730 19818 2790 20435
rect 26237 20408 27037 20438
rect 2957 20362 3023 20365
rect 8845 20362 8911 20365
rect 2957 20360 8911 20362
rect 2957 20304 2962 20360
rect 3018 20304 8850 20360
rect 8906 20304 8911 20360
rect 2957 20302 8911 20304
rect 2957 20299 3023 20302
rect 8845 20299 8911 20302
rect 11697 20362 11763 20365
rect 18873 20362 18939 20365
rect 11697 20360 18939 20362
rect 11697 20304 11702 20360
rect 11758 20304 18878 20360
rect 18934 20304 18939 20360
rect 11697 20302 18939 20304
rect 11697 20299 11763 20302
rect 18873 20299 18939 20302
rect 6821 20226 6887 20229
rect 9213 20226 9279 20229
rect 6821 20224 9279 20226
rect 6821 20168 6826 20224
rect 6882 20168 9218 20224
rect 9274 20168 9279 20224
rect 6821 20166 9279 20168
rect 6821 20163 6887 20166
rect 9213 20163 9279 20166
rect 4039 20160 4355 20161
rect 4039 20096 4045 20160
rect 4109 20096 4125 20160
rect 4189 20096 4205 20160
rect 4269 20096 4285 20160
rect 4349 20096 4355 20160
rect 4039 20095 4355 20096
rect 10226 20160 10542 20161
rect 10226 20096 10232 20160
rect 10296 20096 10312 20160
rect 10376 20096 10392 20160
rect 10456 20096 10472 20160
rect 10536 20096 10542 20160
rect 10226 20095 10542 20096
rect 16413 20160 16729 20161
rect 16413 20096 16419 20160
rect 16483 20096 16499 20160
rect 16563 20096 16579 20160
rect 16643 20096 16659 20160
rect 16723 20096 16729 20160
rect 16413 20095 16729 20096
rect 22600 20160 22916 20161
rect 22600 20096 22606 20160
rect 22670 20096 22686 20160
rect 22750 20096 22766 20160
rect 22830 20096 22846 20160
rect 22910 20096 22916 20160
rect 22600 20095 22916 20096
rect 8477 20090 8543 20093
rect 4478 20088 8543 20090
rect 4478 20032 8482 20088
rect 8538 20032 8543 20088
rect 4478 20030 8543 20032
rect 4245 19954 4311 19957
rect 4478 19954 4538 20030
rect 8477 20027 8543 20030
rect 10685 20090 10751 20093
rect 12985 20090 13051 20093
rect 10685 20088 13051 20090
rect 10685 20032 10690 20088
rect 10746 20032 12990 20088
rect 13046 20032 13051 20088
rect 10685 20030 13051 20032
rect 10685 20027 10751 20030
rect 12985 20027 13051 20030
rect 4245 19952 4538 19954
rect 4245 19896 4250 19952
rect 4306 19896 4538 19952
rect 4245 19894 4538 19896
rect 7281 19954 7347 19957
rect 15101 19954 15167 19957
rect 7281 19952 15167 19954
rect 7281 19896 7286 19952
rect 7342 19896 15106 19952
rect 15162 19896 15167 19952
rect 7281 19894 15167 19896
rect 4245 19891 4311 19894
rect 7281 19891 7347 19894
rect 15101 19891 15167 19894
rect 23841 19818 23907 19821
rect 0 19728 858 19818
rect 2730 19816 23907 19818
rect 2730 19760 23846 19816
rect 23902 19760 23907 19816
rect 2730 19758 23907 19760
rect 23841 19755 23907 19758
rect 25957 19818 26023 19821
rect 26237 19818 27037 19848
rect 25957 19816 27037 19818
rect 25957 19760 25962 19816
rect 26018 19760 27037 19816
rect 25957 19758 27037 19760
rect 25957 19755 26023 19758
rect 26237 19728 27037 19758
rect 798 19546 858 19728
rect 4699 19616 5015 19617
rect 4699 19552 4705 19616
rect 4769 19552 4785 19616
rect 4849 19552 4865 19616
rect 4929 19552 4945 19616
rect 5009 19552 5015 19616
rect 4699 19551 5015 19552
rect 10886 19616 11202 19617
rect 10886 19552 10892 19616
rect 10956 19552 10972 19616
rect 11036 19552 11052 19616
rect 11116 19552 11132 19616
rect 11196 19552 11202 19616
rect 10886 19551 11202 19552
rect 17073 19616 17389 19617
rect 17073 19552 17079 19616
rect 17143 19552 17159 19616
rect 17223 19552 17239 19616
rect 17303 19552 17319 19616
rect 17383 19552 17389 19616
rect 17073 19551 17389 19552
rect 23260 19616 23576 19617
rect 23260 19552 23266 19616
rect 23330 19552 23346 19616
rect 23410 19552 23426 19616
rect 23490 19552 23506 19616
rect 23570 19552 23576 19616
rect 23260 19551 23576 19552
rect 1577 19546 1643 19549
rect 798 19544 1643 19546
rect 798 19488 1582 19544
rect 1638 19488 1643 19544
rect 798 19486 1643 19488
rect 1577 19483 1643 19486
rect 1485 19410 1551 19413
rect 19425 19410 19491 19413
rect 1485 19408 19491 19410
rect 1485 19352 1490 19408
rect 1546 19352 19430 19408
rect 19486 19352 19491 19408
rect 1485 19350 19491 19352
rect 1485 19347 1551 19350
rect 19425 19347 19491 19350
rect 1945 19274 2011 19277
rect 982 19272 2011 19274
rect 982 19216 1950 19272
rect 2006 19216 2011 19272
rect 982 19214 2011 19216
rect 0 19138 800 19168
rect 982 19138 1042 19214
rect 1945 19211 2011 19214
rect 4521 19274 4587 19277
rect 8293 19274 8359 19277
rect 4521 19272 8359 19274
rect 4521 19216 4526 19272
rect 4582 19216 8298 19272
rect 8354 19216 8359 19272
rect 4521 19214 8359 19216
rect 4521 19211 4587 19214
rect 8293 19211 8359 19214
rect 12341 19274 12407 19277
rect 12617 19274 12683 19277
rect 18781 19274 18847 19277
rect 12341 19272 18847 19274
rect 12341 19216 12346 19272
rect 12402 19216 12622 19272
rect 12678 19216 18786 19272
rect 18842 19216 18847 19272
rect 12341 19214 18847 19216
rect 12341 19211 12407 19214
rect 12617 19211 12683 19214
rect 18781 19211 18847 19214
rect 0 19078 1042 19138
rect 25405 19138 25471 19141
rect 26237 19138 27037 19168
rect 25405 19136 27037 19138
rect 25405 19080 25410 19136
rect 25466 19080 27037 19136
rect 25405 19078 27037 19080
rect 0 19048 800 19078
rect 25405 19075 25471 19078
rect 4039 19072 4355 19073
rect 4039 19008 4045 19072
rect 4109 19008 4125 19072
rect 4189 19008 4205 19072
rect 4269 19008 4285 19072
rect 4349 19008 4355 19072
rect 4039 19007 4355 19008
rect 10226 19072 10542 19073
rect 10226 19008 10232 19072
rect 10296 19008 10312 19072
rect 10376 19008 10392 19072
rect 10456 19008 10472 19072
rect 10536 19008 10542 19072
rect 10226 19007 10542 19008
rect 16413 19072 16729 19073
rect 16413 19008 16419 19072
rect 16483 19008 16499 19072
rect 16563 19008 16579 19072
rect 16643 19008 16659 19072
rect 16723 19008 16729 19072
rect 16413 19007 16729 19008
rect 22600 19072 22916 19073
rect 22600 19008 22606 19072
rect 22670 19008 22686 19072
rect 22750 19008 22766 19072
rect 22830 19008 22846 19072
rect 22910 19008 22916 19072
rect 26237 19048 27037 19078
rect 22600 19007 22916 19008
rect 4797 19002 4863 19005
rect 4478 19000 4863 19002
rect 4478 18944 4802 19000
rect 4858 18944 4863 19000
rect 4478 18942 4863 18944
rect 4153 18866 4219 18869
rect 4478 18866 4538 18942
rect 4797 18939 4863 18942
rect 14641 19002 14707 19005
rect 15837 19002 15903 19005
rect 14641 19000 15903 19002
rect 14641 18944 14646 19000
rect 14702 18944 15842 19000
rect 15898 18944 15903 19000
rect 14641 18942 15903 18944
rect 14641 18939 14707 18942
rect 15837 18939 15903 18942
rect 4153 18864 4538 18866
rect 4153 18808 4158 18864
rect 4214 18808 4538 18864
rect 4153 18806 4538 18808
rect 4797 18866 4863 18869
rect 5257 18866 5323 18869
rect 4797 18864 5323 18866
rect 4797 18808 4802 18864
rect 4858 18808 5262 18864
rect 5318 18808 5323 18864
rect 4797 18806 5323 18808
rect 4153 18803 4219 18806
rect 4797 18803 4863 18806
rect 5257 18803 5323 18806
rect 10961 18866 11027 18869
rect 25221 18866 25287 18869
rect 10961 18864 25287 18866
rect 10961 18808 10966 18864
rect 11022 18808 25226 18864
rect 25282 18808 25287 18864
rect 10961 18806 25287 18808
rect 10961 18803 11027 18806
rect 25221 18803 25287 18806
rect 4245 18730 4311 18733
rect 7833 18730 7899 18733
rect 4245 18728 7899 18730
rect 4245 18672 4250 18728
rect 4306 18672 7838 18728
rect 7894 18672 7899 18728
rect 4245 18670 7899 18672
rect 4245 18667 4311 18670
rect 7833 18667 7899 18670
rect 14733 18730 14799 18733
rect 15653 18730 15719 18733
rect 14733 18728 15719 18730
rect 14733 18672 14738 18728
rect 14794 18672 15658 18728
rect 15714 18672 15719 18728
rect 14733 18670 15719 18672
rect 14733 18667 14799 18670
rect 15653 18667 15719 18670
rect 4699 18528 5015 18529
rect 4699 18464 4705 18528
rect 4769 18464 4785 18528
rect 4849 18464 4865 18528
rect 4929 18464 4945 18528
rect 5009 18464 5015 18528
rect 4699 18463 5015 18464
rect 10886 18528 11202 18529
rect 10886 18464 10892 18528
rect 10956 18464 10972 18528
rect 11036 18464 11052 18528
rect 11116 18464 11132 18528
rect 11196 18464 11202 18528
rect 10886 18463 11202 18464
rect 17073 18528 17389 18529
rect 17073 18464 17079 18528
rect 17143 18464 17159 18528
rect 17223 18464 17239 18528
rect 17303 18464 17319 18528
rect 17383 18464 17389 18528
rect 17073 18463 17389 18464
rect 23260 18528 23576 18529
rect 23260 18464 23266 18528
rect 23330 18464 23346 18528
rect 23410 18464 23426 18528
rect 23490 18464 23506 18528
rect 23570 18464 23576 18528
rect 23260 18463 23576 18464
rect 25957 18458 26023 18461
rect 26237 18458 27037 18488
rect 25957 18456 27037 18458
rect 25957 18400 25962 18456
rect 26018 18400 27037 18456
rect 25957 18398 27037 18400
rect 25957 18395 26023 18398
rect 26237 18368 27037 18398
rect 1485 18322 1551 18325
rect 15101 18322 15167 18325
rect 16665 18322 16731 18325
rect 1485 18320 2790 18322
rect 1485 18264 1490 18320
rect 1546 18264 2790 18320
rect 1485 18262 2790 18264
rect 1485 18259 1551 18262
rect 2730 18186 2790 18262
rect 15101 18320 16731 18322
rect 15101 18264 15106 18320
rect 15162 18264 16670 18320
rect 16726 18264 16731 18320
rect 15101 18262 16731 18264
rect 15101 18259 15167 18262
rect 16665 18259 16731 18262
rect 2730 18126 16866 18186
rect 16806 18050 16866 18126
rect 18965 18050 19031 18053
rect 21541 18050 21607 18053
rect 16806 18048 21607 18050
rect 16806 17992 18970 18048
rect 19026 17992 21546 18048
rect 21602 17992 21607 18048
rect 16806 17990 21607 17992
rect 18965 17987 19031 17990
rect 21541 17987 21607 17990
rect 4039 17984 4355 17985
rect 4039 17920 4045 17984
rect 4109 17920 4125 17984
rect 4189 17920 4205 17984
rect 4269 17920 4285 17984
rect 4349 17920 4355 17984
rect 4039 17919 4355 17920
rect 10226 17984 10542 17985
rect 10226 17920 10232 17984
rect 10296 17920 10312 17984
rect 10376 17920 10392 17984
rect 10456 17920 10472 17984
rect 10536 17920 10542 17984
rect 10226 17919 10542 17920
rect 16413 17984 16729 17985
rect 16413 17920 16419 17984
rect 16483 17920 16499 17984
rect 16563 17920 16579 17984
rect 16643 17920 16659 17984
rect 16723 17920 16729 17984
rect 16413 17919 16729 17920
rect 22600 17984 22916 17985
rect 22600 17920 22606 17984
rect 22670 17920 22686 17984
rect 22750 17920 22766 17984
rect 22830 17920 22846 17984
rect 22910 17920 22916 17984
rect 22600 17919 22916 17920
rect 1577 17914 1643 17917
rect 798 17912 1643 17914
rect 798 17856 1582 17912
rect 1638 17856 1643 17912
rect 798 17854 1643 17856
rect 798 17808 858 17854
rect 1577 17851 1643 17854
rect 5257 17914 5323 17917
rect 7782 17914 7788 17916
rect 5257 17912 7788 17914
rect 5257 17856 5262 17912
rect 5318 17856 7788 17912
rect 5257 17854 7788 17856
rect 5257 17851 5323 17854
rect 7782 17852 7788 17854
rect 7852 17852 7858 17916
rect 0 17718 858 17808
rect 5441 17778 5507 17781
rect 9673 17778 9739 17781
rect 5441 17776 9739 17778
rect 5441 17720 5446 17776
rect 5502 17720 9678 17776
rect 9734 17720 9739 17776
rect 5441 17718 9739 17720
rect 0 17688 800 17718
rect 5441 17715 5507 17718
rect 9673 17715 9739 17718
rect 5533 17642 5599 17645
rect 11881 17642 11947 17645
rect 5533 17640 11947 17642
rect 5533 17584 5538 17640
rect 5594 17584 11886 17640
rect 11942 17584 11947 17640
rect 5533 17582 11947 17584
rect 5533 17579 5599 17582
rect 11881 17579 11947 17582
rect 4699 17440 5015 17441
rect 4699 17376 4705 17440
rect 4769 17376 4785 17440
rect 4849 17376 4865 17440
rect 4929 17376 4945 17440
rect 5009 17376 5015 17440
rect 4699 17375 5015 17376
rect 10886 17440 11202 17441
rect 10886 17376 10892 17440
rect 10956 17376 10972 17440
rect 11036 17376 11052 17440
rect 11116 17376 11132 17440
rect 11196 17376 11202 17440
rect 10886 17375 11202 17376
rect 17073 17440 17389 17441
rect 17073 17376 17079 17440
rect 17143 17376 17159 17440
rect 17223 17376 17239 17440
rect 17303 17376 17319 17440
rect 17383 17376 17389 17440
rect 17073 17375 17389 17376
rect 23260 17440 23576 17441
rect 23260 17376 23266 17440
rect 23330 17376 23346 17440
rect 23410 17376 23426 17440
rect 23490 17376 23506 17440
rect 23570 17376 23576 17440
rect 23260 17375 23576 17376
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 1577 17098 1643 17101
rect 19609 17098 19675 17101
rect 1577 17096 19675 17098
rect 1577 17040 1582 17096
rect 1638 17040 19614 17096
rect 19670 17040 19675 17096
rect 1577 17038 19675 17040
rect 1577 17035 1643 17038
rect 19609 17035 19675 17038
rect 25681 17098 25747 17101
rect 26237 17098 27037 17128
rect 25681 17096 27037 17098
rect 25681 17040 25686 17096
rect 25742 17040 27037 17096
rect 25681 17038 27037 17040
rect 25681 17035 25747 17038
rect 26237 17008 27037 17038
rect 4039 16896 4355 16897
rect 4039 16832 4045 16896
rect 4109 16832 4125 16896
rect 4189 16832 4205 16896
rect 4269 16832 4285 16896
rect 4349 16832 4355 16896
rect 4039 16831 4355 16832
rect 10226 16896 10542 16897
rect 10226 16832 10232 16896
rect 10296 16832 10312 16896
rect 10376 16832 10392 16896
rect 10456 16832 10472 16896
rect 10536 16832 10542 16896
rect 10226 16831 10542 16832
rect 16413 16896 16729 16897
rect 16413 16832 16419 16896
rect 16483 16832 16499 16896
rect 16563 16832 16579 16896
rect 16643 16832 16659 16896
rect 16723 16832 16729 16896
rect 16413 16831 16729 16832
rect 22600 16896 22916 16897
rect 22600 16832 22606 16896
rect 22670 16832 22686 16896
rect 22750 16832 22766 16896
rect 22830 16832 22846 16896
rect 22910 16832 22916 16896
rect 22600 16831 22916 16832
rect 13813 16690 13879 16693
rect 18965 16690 19031 16693
rect 13813 16688 19031 16690
rect 13813 16632 13818 16688
rect 13874 16632 18970 16688
rect 19026 16632 19031 16688
rect 13813 16630 19031 16632
rect 13813 16627 13879 16630
rect 18965 16627 19031 16630
rect 1393 16554 1459 16557
rect 798 16552 1459 16554
rect 798 16496 1398 16552
rect 1454 16496 1459 16552
rect 798 16494 1459 16496
rect 798 16448 858 16494
rect 1393 16491 1459 16494
rect 5441 16554 5507 16557
rect 8937 16554 9003 16557
rect 5441 16552 9003 16554
rect 5441 16496 5446 16552
rect 5502 16496 8942 16552
rect 8998 16496 9003 16552
rect 5441 16494 9003 16496
rect 5441 16491 5507 16494
rect 8937 16491 9003 16494
rect 10501 16554 10567 16557
rect 12525 16554 12591 16557
rect 18413 16554 18479 16557
rect 10501 16552 12591 16554
rect 10501 16496 10506 16552
rect 10562 16496 12530 16552
rect 12586 16496 12591 16552
rect 10501 16494 12591 16496
rect 10501 16491 10567 16494
rect 12525 16491 12591 16494
rect 15840 16552 18479 16554
rect 15840 16496 18418 16552
rect 18474 16496 18479 16552
rect 15840 16494 18479 16496
rect 0 16358 858 16448
rect 11421 16418 11487 16421
rect 15840 16418 15900 16494
rect 18413 16491 18479 16494
rect 11421 16416 15900 16418
rect 11421 16360 11426 16416
rect 11482 16360 15900 16416
rect 11421 16358 15900 16360
rect 25957 16418 26023 16421
rect 26237 16418 27037 16448
rect 25957 16416 27037 16418
rect 25957 16360 25962 16416
rect 26018 16360 27037 16416
rect 25957 16358 27037 16360
rect 0 16328 800 16358
rect 11421 16355 11487 16358
rect 25957 16355 26023 16358
rect 4699 16352 5015 16353
rect 4699 16288 4705 16352
rect 4769 16288 4785 16352
rect 4849 16288 4865 16352
rect 4929 16288 4945 16352
rect 5009 16288 5015 16352
rect 4699 16287 5015 16288
rect 10886 16352 11202 16353
rect 10886 16288 10892 16352
rect 10956 16288 10972 16352
rect 11036 16288 11052 16352
rect 11116 16288 11132 16352
rect 11196 16288 11202 16352
rect 10886 16287 11202 16288
rect 17073 16352 17389 16353
rect 17073 16288 17079 16352
rect 17143 16288 17159 16352
rect 17223 16288 17239 16352
rect 17303 16288 17319 16352
rect 17383 16288 17389 16352
rect 17073 16287 17389 16288
rect 23260 16352 23576 16353
rect 23260 16288 23266 16352
rect 23330 16288 23346 16352
rect 23410 16288 23426 16352
rect 23490 16288 23506 16352
rect 23570 16288 23576 16352
rect 26237 16328 27037 16358
rect 23260 16287 23576 16288
rect 1853 16146 1919 16149
rect 23197 16146 23263 16149
rect 1853 16144 23263 16146
rect 1853 16088 1858 16144
rect 1914 16088 23202 16144
rect 23258 16088 23263 16144
rect 1853 16086 23263 16088
rect 1853 16083 1919 16086
rect 23197 16083 23263 16086
rect 23381 16146 23447 16149
rect 25037 16146 25103 16149
rect 23381 16144 25103 16146
rect 23381 16088 23386 16144
rect 23442 16088 25042 16144
rect 25098 16088 25103 16144
rect 23381 16086 25103 16088
rect 23381 16083 23447 16086
rect 25037 16083 25103 16086
rect 11237 16010 11303 16013
rect 22369 16010 22435 16013
rect 11237 16008 22435 16010
rect 11237 15952 11242 16008
rect 11298 15952 22374 16008
rect 22430 15952 22435 16008
rect 11237 15950 22435 15952
rect 11237 15947 11303 15950
rect 22369 15947 22435 15950
rect 4039 15808 4355 15809
rect 0 15738 800 15768
rect 4039 15744 4045 15808
rect 4109 15744 4125 15808
rect 4189 15744 4205 15808
rect 4269 15744 4285 15808
rect 4349 15744 4355 15808
rect 4039 15743 4355 15744
rect 10226 15808 10542 15809
rect 10226 15744 10232 15808
rect 10296 15744 10312 15808
rect 10376 15744 10392 15808
rect 10456 15744 10472 15808
rect 10536 15744 10542 15808
rect 10226 15743 10542 15744
rect 16413 15808 16729 15809
rect 16413 15744 16419 15808
rect 16483 15744 16499 15808
rect 16563 15744 16579 15808
rect 16643 15744 16659 15808
rect 16723 15744 16729 15808
rect 16413 15743 16729 15744
rect 22600 15808 22916 15809
rect 22600 15744 22606 15808
rect 22670 15744 22686 15808
rect 22750 15744 22766 15808
rect 22830 15744 22846 15808
rect 22910 15744 22916 15808
rect 22600 15743 22916 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 25405 15738 25471 15741
rect 26237 15738 27037 15768
rect 25405 15736 27037 15738
rect 25405 15680 25410 15736
rect 25466 15680 27037 15736
rect 25405 15678 27037 15680
rect 25405 15675 25471 15678
rect 26237 15648 27037 15678
rect 1761 15466 1827 15469
rect 23933 15466 23999 15469
rect 1761 15464 23999 15466
rect 1761 15408 1766 15464
rect 1822 15408 23938 15464
rect 23994 15408 23999 15464
rect 1761 15406 23999 15408
rect 1761 15403 1827 15406
rect 23933 15403 23999 15406
rect 4699 15264 5015 15265
rect 4699 15200 4705 15264
rect 4769 15200 4785 15264
rect 4849 15200 4865 15264
rect 4929 15200 4945 15264
rect 5009 15200 5015 15264
rect 4699 15199 5015 15200
rect 10886 15264 11202 15265
rect 10886 15200 10892 15264
rect 10956 15200 10972 15264
rect 11036 15200 11052 15264
rect 11116 15200 11132 15264
rect 11196 15200 11202 15264
rect 10886 15199 11202 15200
rect 17073 15264 17389 15265
rect 17073 15200 17079 15264
rect 17143 15200 17159 15264
rect 17223 15200 17239 15264
rect 17303 15200 17319 15264
rect 17383 15200 17389 15264
rect 17073 15199 17389 15200
rect 23260 15264 23576 15265
rect 23260 15200 23266 15264
rect 23330 15200 23346 15264
rect 23410 15200 23426 15264
rect 23490 15200 23506 15264
rect 23570 15200 23576 15264
rect 23260 15199 23576 15200
rect 8845 15058 8911 15061
rect 15193 15058 15259 15061
rect 8845 15056 15259 15058
rect 8845 15000 8850 15056
rect 8906 15000 15198 15056
rect 15254 15000 15259 15056
rect 8845 14998 15259 15000
rect 8845 14995 8911 14998
rect 15193 14995 15259 14998
rect 4039 14720 4355 14721
rect 4039 14656 4045 14720
rect 4109 14656 4125 14720
rect 4189 14656 4205 14720
rect 4269 14656 4285 14720
rect 4349 14656 4355 14720
rect 4039 14655 4355 14656
rect 10226 14720 10542 14721
rect 10226 14656 10232 14720
rect 10296 14656 10312 14720
rect 10376 14656 10392 14720
rect 10456 14656 10472 14720
rect 10536 14656 10542 14720
rect 10226 14655 10542 14656
rect 16413 14720 16729 14721
rect 16413 14656 16419 14720
rect 16483 14656 16499 14720
rect 16563 14656 16579 14720
rect 16643 14656 16659 14720
rect 16723 14656 16729 14720
rect 16413 14655 16729 14656
rect 22600 14720 22916 14721
rect 22600 14656 22606 14720
rect 22670 14656 22686 14720
rect 22750 14656 22766 14720
rect 22830 14656 22846 14720
rect 22910 14656 22916 14720
rect 22600 14655 22916 14656
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 13997 14378 14063 14381
rect 22185 14378 22251 14381
rect 13997 14376 22251 14378
rect 13997 14320 14002 14376
rect 14058 14320 22190 14376
rect 22246 14320 22251 14376
rect 13997 14318 22251 14320
rect 13997 14315 14063 14318
rect 22185 14315 22251 14318
rect 25957 14378 26023 14381
rect 26237 14378 27037 14408
rect 25957 14376 27037 14378
rect 25957 14320 25962 14376
rect 26018 14320 27037 14376
rect 25957 14318 27037 14320
rect 25957 14315 26023 14318
rect 26237 14288 27037 14318
rect 4699 14176 5015 14177
rect 4699 14112 4705 14176
rect 4769 14112 4785 14176
rect 4849 14112 4865 14176
rect 4929 14112 4945 14176
rect 5009 14112 5015 14176
rect 4699 14111 5015 14112
rect 10886 14176 11202 14177
rect 10886 14112 10892 14176
rect 10956 14112 10972 14176
rect 11036 14112 11052 14176
rect 11116 14112 11132 14176
rect 11196 14112 11202 14176
rect 10886 14111 11202 14112
rect 17073 14176 17389 14177
rect 17073 14112 17079 14176
rect 17143 14112 17159 14176
rect 17223 14112 17239 14176
rect 17303 14112 17319 14176
rect 17383 14112 17389 14176
rect 17073 14111 17389 14112
rect 23260 14176 23576 14177
rect 23260 14112 23266 14176
rect 23330 14112 23346 14176
rect 23410 14112 23426 14176
rect 23490 14112 23506 14176
rect 23570 14112 23576 14176
rect 23260 14111 23576 14112
rect 10501 13834 10567 13837
rect 10777 13834 10843 13837
rect 10501 13832 10843 13834
rect 10501 13776 10506 13832
rect 10562 13776 10782 13832
rect 10838 13776 10843 13832
rect 10501 13774 10843 13776
rect 10501 13771 10567 13774
rect 10777 13771 10843 13774
rect 11513 13834 11579 13837
rect 12065 13834 12131 13837
rect 11513 13832 12131 13834
rect 11513 13776 11518 13832
rect 11574 13776 12070 13832
rect 12126 13776 12131 13832
rect 11513 13774 12131 13776
rect 11513 13771 11579 13774
rect 12065 13771 12131 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 25681 13698 25747 13701
rect 26237 13698 27037 13728
rect 25681 13696 27037 13698
rect 25681 13640 25686 13696
rect 25742 13640 27037 13696
rect 25681 13638 27037 13640
rect 25681 13635 25747 13638
rect 4039 13632 4355 13633
rect 4039 13568 4045 13632
rect 4109 13568 4125 13632
rect 4189 13568 4205 13632
rect 4269 13568 4285 13632
rect 4349 13568 4355 13632
rect 4039 13567 4355 13568
rect 10226 13632 10542 13633
rect 10226 13568 10232 13632
rect 10296 13568 10312 13632
rect 10376 13568 10392 13632
rect 10456 13568 10472 13632
rect 10536 13568 10542 13632
rect 10226 13567 10542 13568
rect 16413 13632 16729 13633
rect 16413 13568 16419 13632
rect 16483 13568 16499 13632
rect 16563 13568 16579 13632
rect 16643 13568 16659 13632
rect 16723 13568 16729 13632
rect 16413 13567 16729 13568
rect 22600 13632 22916 13633
rect 22600 13568 22606 13632
rect 22670 13568 22686 13632
rect 22750 13568 22766 13632
rect 22830 13568 22846 13632
rect 22910 13568 22916 13632
rect 26237 13608 27037 13638
rect 22600 13567 22916 13568
rect 6453 13426 6519 13429
rect 16573 13426 16639 13429
rect 6453 13424 16639 13426
rect 6453 13368 6458 13424
rect 6514 13368 16578 13424
rect 16634 13368 16639 13424
rect 6453 13366 16639 13368
rect 6453 13363 6519 13366
rect 16573 13363 16639 13366
rect 4337 13290 4403 13293
rect 8109 13290 8175 13293
rect 4337 13288 8175 13290
rect 4337 13232 4342 13288
rect 4398 13232 8114 13288
rect 8170 13232 8175 13288
rect 4337 13230 8175 13232
rect 4337 13227 4403 13230
rect 8109 13227 8175 13230
rect 9765 13290 9831 13293
rect 20529 13290 20595 13293
rect 9765 13288 20595 13290
rect 9765 13232 9770 13288
rect 9826 13232 20534 13288
rect 20590 13232 20595 13288
rect 9765 13230 20595 13232
rect 9765 13227 9831 13230
rect 20529 13227 20595 13230
rect 4699 13088 5015 13089
rect 0 13018 800 13048
rect 4699 13024 4705 13088
rect 4769 13024 4785 13088
rect 4849 13024 4865 13088
rect 4929 13024 4945 13088
rect 5009 13024 5015 13088
rect 4699 13023 5015 13024
rect 10886 13088 11202 13089
rect 10886 13024 10892 13088
rect 10956 13024 10972 13088
rect 11036 13024 11052 13088
rect 11116 13024 11132 13088
rect 11196 13024 11202 13088
rect 10886 13023 11202 13024
rect 17073 13088 17389 13089
rect 17073 13024 17079 13088
rect 17143 13024 17159 13088
rect 17223 13024 17239 13088
rect 17303 13024 17319 13088
rect 17383 13024 17389 13088
rect 17073 13023 17389 13024
rect 23260 13088 23576 13089
rect 23260 13024 23266 13088
rect 23330 13024 23346 13088
rect 23410 13024 23426 13088
rect 23490 13024 23506 13088
rect 23570 13024 23576 13088
rect 23260 13023 23576 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 25405 13018 25471 13021
rect 26237 13018 27037 13048
rect 25405 13016 27037 13018
rect 25405 12960 25410 13016
rect 25466 12960 27037 13016
rect 25405 12958 27037 12960
rect 25405 12955 25471 12958
rect 26237 12928 27037 12958
rect 11881 12882 11947 12885
rect 11881 12880 22110 12882
rect 11881 12824 11886 12880
rect 11942 12824 22110 12880
rect 11881 12822 22110 12824
rect 11881 12819 11947 12822
rect 12709 12746 12775 12749
rect 15837 12746 15903 12749
rect 12709 12744 15903 12746
rect 12709 12688 12714 12744
rect 12770 12688 15842 12744
rect 15898 12688 15903 12744
rect 12709 12686 15903 12688
rect 22050 12746 22110 12822
rect 26325 12746 26391 12749
rect 22050 12744 26391 12746
rect 22050 12688 26330 12744
rect 26386 12688 26391 12744
rect 22050 12686 26391 12688
rect 12709 12683 12775 12686
rect 15837 12683 15903 12686
rect 26325 12683 26391 12686
rect 4039 12544 4355 12545
rect 4039 12480 4045 12544
rect 4109 12480 4125 12544
rect 4189 12480 4205 12544
rect 4269 12480 4285 12544
rect 4349 12480 4355 12544
rect 4039 12479 4355 12480
rect 10226 12544 10542 12545
rect 10226 12480 10232 12544
rect 10296 12480 10312 12544
rect 10376 12480 10392 12544
rect 10456 12480 10472 12544
rect 10536 12480 10542 12544
rect 10226 12479 10542 12480
rect 16413 12544 16729 12545
rect 16413 12480 16419 12544
rect 16483 12480 16499 12544
rect 16563 12480 16579 12544
rect 16643 12480 16659 12544
rect 16723 12480 16729 12544
rect 16413 12479 16729 12480
rect 22600 12544 22916 12545
rect 22600 12480 22606 12544
rect 22670 12480 22686 12544
rect 22750 12480 22766 12544
rect 22830 12480 22846 12544
rect 22910 12480 22916 12544
rect 22600 12479 22916 12480
rect 11053 12338 11119 12341
rect 11881 12338 11947 12341
rect 11053 12336 11947 12338
rect 11053 12280 11058 12336
rect 11114 12280 11886 12336
rect 11942 12280 11947 12336
rect 11053 12278 11947 12280
rect 11053 12275 11119 12278
rect 11881 12275 11947 12278
rect 26049 12338 26115 12341
rect 26237 12338 27037 12368
rect 26049 12336 27037 12338
rect 26049 12280 26054 12336
rect 26110 12280 27037 12336
rect 26049 12278 27037 12280
rect 26049 12275 26115 12278
rect 26237 12248 27037 12278
rect 6085 12202 6151 12205
rect 11973 12202 12039 12205
rect 6085 12200 12039 12202
rect 6085 12144 6090 12200
rect 6146 12144 11978 12200
rect 12034 12144 12039 12200
rect 6085 12142 12039 12144
rect 6085 12139 6151 12142
rect 11973 12139 12039 12142
rect 4699 12000 5015 12001
rect 4699 11936 4705 12000
rect 4769 11936 4785 12000
rect 4849 11936 4865 12000
rect 4929 11936 4945 12000
rect 5009 11936 5015 12000
rect 4699 11935 5015 11936
rect 10886 12000 11202 12001
rect 10886 11936 10892 12000
rect 10956 11936 10972 12000
rect 11036 11936 11052 12000
rect 11116 11936 11132 12000
rect 11196 11936 11202 12000
rect 10886 11935 11202 11936
rect 17073 12000 17389 12001
rect 17073 11936 17079 12000
rect 17143 11936 17159 12000
rect 17223 11936 17239 12000
rect 17303 11936 17319 12000
rect 17383 11936 17389 12000
rect 17073 11935 17389 11936
rect 23260 12000 23576 12001
rect 23260 11936 23266 12000
rect 23330 11936 23346 12000
rect 23410 11936 23426 12000
rect 23490 11936 23506 12000
rect 23570 11936 23576 12000
rect 23260 11935 23576 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 15326 11596 15332 11660
rect 15396 11658 15402 11660
rect 15837 11658 15903 11661
rect 15396 11656 15903 11658
rect 15396 11600 15842 11656
rect 15898 11600 15903 11656
rect 15396 11598 15903 11600
rect 15396 11596 15402 11598
rect 15837 11595 15903 11598
rect 4039 11456 4355 11457
rect 4039 11392 4045 11456
rect 4109 11392 4125 11456
rect 4189 11392 4205 11456
rect 4269 11392 4285 11456
rect 4349 11392 4355 11456
rect 4039 11391 4355 11392
rect 10226 11456 10542 11457
rect 10226 11392 10232 11456
rect 10296 11392 10312 11456
rect 10376 11392 10392 11456
rect 10456 11392 10472 11456
rect 10536 11392 10542 11456
rect 10226 11391 10542 11392
rect 16413 11456 16729 11457
rect 16413 11392 16419 11456
rect 16483 11392 16499 11456
rect 16563 11392 16579 11456
rect 16643 11392 16659 11456
rect 16723 11392 16729 11456
rect 16413 11391 16729 11392
rect 22600 11456 22916 11457
rect 22600 11392 22606 11456
rect 22670 11392 22686 11456
rect 22750 11392 22766 11456
rect 22830 11392 22846 11456
rect 22910 11392 22916 11456
rect 22600 11391 22916 11392
rect 13905 11114 13971 11117
rect 17309 11114 17375 11117
rect 13905 11112 17375 11114
rect 13905 11056 13910 11112
rect 13966 11056 17314 11112
rect 17370 11056 17375 11112
rect 13905 11054 17375 11056
rect 13905 11051 13971 11054
rect 17309 11051 17375 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 25957 10978 26023 10981
rect 26237 10978 27037 11008
rect 25957 10976 27037 10978
rect 25957 10920 25962 10976
rect 26018 10920 27037 10976
rect 25957 10918 27037 10920
rect 25957 10915 26023 10918
rect 4699 10912 5015 10913
rect 4699 10848 4705 10912
rect 4769 10848 4785 10912
rect 4849 10848 4865 10912
rect 4929 10848 4945 10912
rect 5009 10848 5015 10912
rect 4699 10847 5015 10848
rect 10886 10912 11202 10913
rect 10886 10848 10892 10912
rect 10956 10848 10972 10912
rect 11036 10848 11052 10912
rect 11116 10848 11132 10912
rect 11196 10848 11202 10912
rect 10886 10847 11202 10848
rect 17073 10912 17389 10913
rect 17073 10848 17079 10912
rect 17143 10848 17159 10912
rect 17223 10848 17239 10912
rect 17303 10848 17319 10912
rect 17383 10848 17389 10912
rect 17073 10847 17389 10848
rect 23260 10912 23576 10913
rect 23260 10848 23266 10912
rect 23330 10848 23346 10912
rect 23410 10848 23426 10912
rect 23490 10848 23506 10912
rect 23570 10848 23576 10912
rect 26237 10888 27037 10918
rect 23260 10847 23576 10848
rect 1485 10706 1551 10709
rect 20713 10706 20779 10709
rect 1485 10704 20779 10706
rect 1485 10648 1490 10704
rect 1546 10648 20718 10704
rect 20774 10648 20779 10704
rect 1485 10646 20779 10648
rect 1485 10643 1551 10646
rect 20713 10643 20779 10646
rect 5073 10570 5139 10573
rect 5533 10570 5599 10573
rect 17125 10570 17191 10573
rect 5073 10568 5599 10570
rect 5073 10512 5078 10568
rect 5134 10512 5538 10568
rect 5594 10512 5599 10568
rect 5073 10510 5599 10512
rect 5073 10507 5139 10510
rect 5533 10507 5599 10510
rect 16254 10568 17191 10570
rect 16254 10512 17130 10568
rect 17186 10512 17191 10568
rect 16254 10510 17191 10512
rect 4039 10368 4355 10369
rect 0 10298 800 10328
rect 4039 10304 4045 10368
rect 4109 10304 4125 10368
rect 4189 10304 4205 10368
rect 4269 10304 4285 10368
rect 4349 10304 4355 10368
rect 4039 10303 4355 10304
rect 10226 10368 10542 10369
rect 10226 10304 10232 10368
rect 10296 10304 10312 10368
rect 10376 10304 10392 10368
rect 10456 10304 10472 10368
rect 10536 10304 10542 10368
rect 10226 10303 10542 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 12893 10298 12959 10301
rect 14825 10298 14891 10301
rect 16254 10298 16314 10510
rect 17125 10507 17191 10510
rect 16413 10368 16729 10369
rect 16413 10304 16419 10368
rect 16483 10304 16499 10368
rect 16563 10304 16579 10368
rect 16643 10304 16659 10368
rect 16723 10304 16729 10368
rect 16413 10303 16729 10304
rect 22600 10368 22916 10369
rect 22600 10304 22606 10368
rect 22670 10304 22686 10368
rect 22750 10304 22766 10368
rect 22830 10304 22846 10368
rect 22910 10304 22916 10368
rect 22600 10303 22916 10304
rect 12893 10296 16314 10298
rect 12893 10240 12898 10296
rect 12954 10240 14830 10296
rect 14886 10240 16314 10296
rect 12893 10238 16314 10240
rect 25405 10298 25471 10301
rect 26237 10298 27037 10328
rect 25405 10296 27037 10298
rect 25405 10240 25410 10296
rect 25466 10240 27037 10296
rect 25405 10238 27037 10240
rect 12893 10235 12959 10238
rect 14825 10235 14891 10238
rect 25405 10235 25471 10238
rect 26237 10208 27037 10238
rect 1669 10162 1735 10165
rect 19609 10162 19675 10165
rect 1669 10160 19675 10162
rect 1669 10104 1674 10160
rect 1730 10104 19614 10160
rect 19670 10104 19675 10160
rect 1669 10102 19675 10104
rect 1669 10099 1735 10102
rect 19609 10099 19675 10102
rect 2129 10026 2195 10029
rect 24945 10026 25011 10029
rect 2129 10024 25011 10026
rect 2129 9968 2134 10024
rect 2190 9968 24950 10024
rect 25006 9968 25011 10024
rect 2129 9966 25011 9968
rect 2129 9963 2195 9966
rect 24945 9963 25011 9966
rect 12525 9890 12591 9893
rect 16573 9890 16639 9893
rect 16941 9890 17007 9893
rect 17769 9890 17835 9893
rect 12525 9888 16639 9890
rect 12525 9832 12530 9888
rect 12586 9832 16578 9888
rect 16634 9832 16639 9888
rect 12525 9830 16639 9832
rect 12525 9827 12591 9830
rect 16573 9827 16639 9830
rect 16806 9888 17007 9890
rect 16806 9832 16946 9888
rect 17002 9832 17007 9888
rect 16806 9830 17007 9832
rect 4699 9824 5015 9825
rect 4699 9760 4705 9824
rect 4769 9760 4785 9824
rect 4849 9760 4865 9824
rect 4929 9760 4945 9824
rect 5009 9760 5015 9824
rect 4699 9759 5015 9760
rect 10886 9824 11202 9825
rect 10886 9760 10892 9824
rect 10956 9760 10972 9824
rect 11036 9760 11052 9824
rect 11116 9760 11132 9824
rect 11196 9760 11202 9824
rect 10886 9759 11202 9760
rect 12525 9754 12591 9757
rect 13261 9754 13327 9757
rect 12525 9752 13327 9754
rect 12525 9696 12530 9752
rect 12586 9696 13266 9752
rect 13322 9696 13327 9752
rect 12525 9694 13327 9696
rect 12525 9691 12591 9694
rect 13261 9691 13327 9694
rect 16389 9754 16455 9757
rect 16665 9754 16731 9757
rect 16389 9752 16731 9754
rect 16389 9696 16394 9752
rect 16450 9696 16670 9752
rect 16726 9696 16731 9752
rect 16389 9694 16731 9696
rect 16389 9691 16455 9694
rect 16665 9691 16731 9694
rect 16806 9690 16866 9830
rect 16941 9827 17007 9830
rect 17726 9888 17835 9890
rect 17726 9832 17774 9888
rect 17830 9832 17835 9888
rect 17726 9827 17835 9832
rect 17073 9824 17389 9825
rect 17073 9760 17079 9824
rect 17143 9760 17159 9824
rect 17223 9760 17239 9824
rect 17303 9760 17319 9824
rect 17383 9760 17389 9824
rect 17073 9759 17389 9760
rect 17726 9693 17786 9827
rect 23260 9824 23576 9825
rect 23260 9760 23266 9824
rect 23330 9760 23346 9824
rect 23410 9760 23426 9824
rect 23490 9760 23506 9824
rect 23570 9760 23576 9824
rect 23260 9759 23576 9760
rect 17033 9690 17099 9693
rect 16806 9688 17099 9690
rect 0 9618 800 9648
rect 16806 9632 17038 9688
rect 17094 9632 17099 9688
rect 16806 9630 17099 9632
rect 17033 9627 17099 9630
rect 17677 9688 17786 9693
rect 17677 9632 17682 9688
rect 17738 9632 17786 9688
rect 17677 9630 17786 9632
rect 17677 9627 17743 9630
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 800 9558
rect 933 9555 999 9558
rect 4245 9618 4311 9621
rect 5809 9618 5875 9621
rect 4245 9616 5875 9618
rect 4245 9560 4250 9616
rect 4306 9560 5814 9616
rect 5870 9560 5875 9616
rect 4245 9558 5875 9560
rect 4245 9555 4311 9558
rect 5809 9555 5875 9558
rect 11053 9618 11119 9621
rect 13169 9618 13235 9621
rect 11053 9616 13235 9618
rect 11053 9560 11058 9616
rect 11114 9560 13174 9616
rect 13230 9560 13235 9616
rect 11053 9558 13235 9560
rect 11053 9555 11119 9558
rect 13169 9555 13235 9558
rect 25957 9618 26023 9621
rect 26237 9618 27037 9648
rect 25957 9616 27037 9618
rect 25957 9560 25962 9616
rect 26018 9560 27037 9616
rect 25957 9558 27037 9560
rect 25957 9555 26023 9558
rect 26237 9528 27037 9558
rect 9765 9482 9831 9485
rect 11605 9482 11671 9485
rect 9765 9480 11671 9482
rect 9765 9424 9770 9480
rect 9826 9424 11610 9480
rect 11666 9424 11671 9480
rect 9765 9422 11671 9424
rect 9765 9419 9831 9422
rect 11605 9419 11671 9422
rect 12617 9482 12683 9485
rect 13445 9482 13511 9485
rect 12617 9480 13511 9482
rect 12617 9424 12622 9480
rect 12678 9424 13450 9480
rect 13506 9424 13511 9480
rect 12617 9422 13511 9424
rect 12617 9419 12683 9422
rect 13445 9419 13511 9422
rect 10777 9346 10843 9349
rect 14273 9346 14339 9349
rect 10777 9344 14339 9346
rect 10777 9288 10782 9344
rect 10838 9288 14278 9344
rect 14334 9288 14339 9344
rect 10777 9286 14339 9288
rect 10777 9283 10843 9286
rect 14273 9283 14339 9286
rect 4039 9280 4355 9281
rect 4039 9216 4045 9280
rect 4109 9216 4125 9280
rect 4189 9216 4205 9280
rect 4269 9216 4285 9280
rect 4349 9216 4355 9280
rect 4039 9215 4355 9216
rect 10226 9280 10542 9281
rect 10226 9216 10232 9280
rect 10296 9216 10312 9280
rect 10376 9216 10392 9280
rect 10456 9216 10472 9280
rect 10536 9216 10542 9280
rect 10226 9215 10542 9216
rect 16413 9280 16729 9281
rect 16413 9216 16419 9280
rect 16483 9216 16499 9280
rect 16563 9216 16579 9280
rect 16643 9216 16659 9280
rect 16723 9216 16729 9280
rect 16413 9215 16729 9216
rect 22600 9280 22916 9281
rect 22600 9216 22606 9280
rect 22670 9216 22686 9280
rect 22750 9216 22766 9280
rect 22830 9216 22846 9280
rect 22910 9216 22916 9280
rect 22600 9215 22916 9216
rect 9673 9210 9739 9213
rect 9630 9208 9739 9210
rect 9630 9152 9678 9208
rect 9734 9152 9739 9208
rect 9630 9147 9739 9152
rect 11881 9210 11947 9213
rect 13537 9210 13603 9213
rect 11881 9208 13603 9210
rect 11881 9152 11886 9208
rect 11942 9152 13542 9208
rect 13598 9152 13603 9208
rect 11881 9150 13603 9152
rect 11881 9147 11947 9150
rect 13537 9147 13603 9150
rect 9630 8941 9690 9147
rect 9857 9074 9923 9077
rect 10133 9074 10199 9077
rect 9857 9072 10199 9074
rect 9857 9016 9862 9072
rect 9918 9016 10138 9072
rect 10194 9016 10199 9072
rect 9857 9014 10199 9016
rect 9857 9011 9923 9014
rect 10133 9011 10199 9014
rect 11237 9074 11303 9077
rect 13537 9074 13603 9077
rect 11237 9072 13603 9074
rect 11237 9016 11242 9072
rect 11298 9016 13542 9072
rect 13598 9016 13603 9072
rect 11237 9014 13603 9016
rect 11237 9011 11303 9014
rect 13537 9011 13603 9014
rect 9630 8936 9739 8941
rect 9630 8880 9678 8936
rect 9734 8880 9739 8936
rect 9630 8878 9739 8880
rect 9673 8875 9739 8878
rect 11881 8802 11947 8805
rect 12249 8802 12315 8805
rect 11881 8800 12315 8802
rect 11881 8744 11886 8800
rect 11942 8744 12254 8800
rect 12310 8744 12315 8800
rect 11881 8742 12315 8744
rect 11881 8739 11947 8742
rect 12249 8739 12315 8742
rect 4699 8736 5015 8737
rect 4699 8672 4705 8736
rect 4769 8672 4785 8736
rect 4849 8672 4865 8736
rect 4929 8672 4945 8736
rect 5009 8672 5015 8736
rect 4699 8671 5015 8672
rect 10886 8736 11202 8737
rect 10886 8672 10892 8736
rect 10956 8672 10972 8736
rect 11036 8672 11052 8736
rect 11116 8672 11132 8736
rect 11196 8672 11202 8736
rect 10886 8671 11202 8672
rect 17073 8736 17389 8737
rect 17073 8672 17079 8736
rect 17143 8672 17159 8736
rect 17223 8672 17239 8736
rect 17303 8672 17319 8736
rect 17383 8672 17389 8736
rect 17073 8671 17389 8672
rect 23260 8736 23576 8737
rect 23260 8672 23266 8736
rect 23330 8672 23346 8736
rect 23410 8672 23426 8736
rect 23490 8672 23506 8736
rect 23570 8672 23576 8736
rect 23260 8671 23576 8672
rect 0 8258 800 8288
rect 1669 8258 1735 8261
rect 0 8256 1735 8258
rect 0 8200 1674 8256
rect 1730 8200 1735 8256
rect 0 8198 1735 8200
rect 0 8168 800 8198
rect 1669 8195 1735 8198
rect 25957 8258 26023 8261
rect 26237 8258 27037 8288
rect 25957 8256 27037 8258
rect 25957 8200 25962 8256
rect 26018 8200 27037 8256
rect 25957 8198 27037 8200
rect 25957 8195 26023 8198
rect 4039 8192 4355 8193
rect 4039 8128 4045 8192
rect 4109 8128 4125 8192
rect 4189 8128 4205 8192
rect 4269 8128 4285 8192
rect 4349 8128 4355 8192
rect 4039 8127 4355 8128
rect 10226 8192 10542 8193
rect 10226 8128 10232 8192
rect 10296 8128 10312 8192
rect 10376 8128 10392 8192
rect 10456 8128 10472 8192
rect 10536 8128 10542 8192
rect 10226 8127 10542 8128
rect 16413 8192 16729 8193
rect 16413 8128 16419 8192
rect 16483 8128 16499 8192
rect 16563 8128 16579 8192
rect 16643 8128 16659 8192
rect 16723 8128 16729 8192
rect 16413 8127 16729 8128
rect 22600 8192 22916 8193
rect 22600 8128 22606 8192
rect 22670 8128 22686 8192
rect 22750 8128 22766 8192
rect 22830 8128 22846 8192
rect 22910 8128 22916 8192
rect 26237 8168 27037 8198
rect 22600 8127 22916 8128
rect 6545 7850 6611 7853
rect 7649 7850 7715 7853
rect 6545 7848 7715 7850
rect 6545 7792 6550 7848
rect 6606 7792 7654 7848
rect 7710 7792 7715 7848
rect 6545 7790 7715 7792
rect 6545 7787 6611 7790
rect 7649 7787 7715 7790
rect 4699 7648 5015 7649
rect 0 7578 800 7608
rect 4699 7584 4705 7648
rect 4769 7584 4785 7648
rect 4849 7584 4865 7648
rect 4929 7584 4945 7648
rect 5009 7584 5015 7648
rect 4699 7583 5015 7584
rect 10886 7648 11202 7649
rect 10886 7584 10892 7648
rect 10956 7584 10972 7648
rect 11036 7584 11052 7648
rect 11116 7584 11132 7648
rect 11196 7584 11202 7648
rect 10886 7583 11202 7584
rect 17073 7648 17389 7649
rect 17073 7584 17079 7648
rect 17143 7584 17159 7648
rect 17223 7584 17239 7648
rect 17303 7584 17319 7648
rect 17383 7584 17389 7648
rect 17073 7583 17389 7584
rect 23260 7648 23576 7649
rect 23260 7584 23266 7648
rect 23330 7584 23346 7648
rect 23410 7584 23426 7648
rect 23490 7584 23506 7648
rect 23570 7584 23576 7648
rect 23260 7583 23576 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 25681 7578 25747 7581
rect 26237 7578 27037 7608
rect 25681 7576 27037 7578
rect 25681 7520 25686 7576
rect 25742 7520 27037 7576
rect 25681 7518 27037 7520
rect 25681 7515 25747 7518
rect 26237 7488 27037 7518
rect 17677 7306 17743 7309
rect 17677 7304 17786 7306
rect 17677 7248 17682 7304
rect 17738 7248 17786 7304
rect 17677 7243 17786 7248
rect 7833 7170 7899 7173
rect 8201 7170 8267 7173
rect 7833 7168 8267 7170
rect 7833 7112 7838 7168
rect 7894 7112 8206 7168
rect 8262 7112 8267 7168
rect 7833 7110 8267 7112
rect 7833 7107 7899 7110
rect 8201 7107 8267 7110
rect 4039 7104 4355 7105
rect 4039 7040 4045 7104
rect 4109 7040 4125 7104
rect 4189 7040 4205 7104
rect 4269 7040 4285 7104
rect 4349 7040 4355 7104
rect 4039 7039 4355 7040
rect 10226 7104 10542 7105
rect 10226 7040 10232 7104
rect 10296 7040 10312 7104
rect 10376 7040 10392 7104
rect 10456 7040 10472 7104
rect 10536 7040 10542 7104
rect 10226 7039 10542 7040
rect 16413 7104 16729 7105
rect 16413 7040 16419 7104
rect 16483 7040 16499 7104
rect 16563 7040 16579 7104
rect 16643 7040 16659 7104
rect 16723 7040 16729 7104
rect 16413 7039 16729 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 5349 6762 5415 6765
rect 9581 6762 9647 6765
rect 5349 6760 9647 6762
rect 5349 6704 5354 6760
rect 5410 6704 9586 6760
rect 9642 6704 9647 6760
rect 5349 6702 9647 6704
rect 5349 6699 5415 6702
rect 9581 6699 9647 6702
rect 17726 6629 17786 7243
rect 22600 7104 22916 7105
rect 22600 7040 22606 7104
rect 22670 7040 22686 7104
rect 22750 7040 22766 7104
rect 22830 7040 22846 7104
rect 22910 7040 22916 7104
rect 22600 7039 22916 7040
rect 25957 6898 26023 6901
rect 26237 6898 27037 6928
rect 25957 6896 27037 6898
rect 25957 6840 25962 6896
rect 26018 6840 27037 6896
rect 25957 6838 27037 6840
rect 25957 6835 26023 6838
rect 26237 6808 27037 6838
rect 17726 6624 17835 6629
rect 17726 6568 17774 6624
rect 17830 6568 17835 6624
rect 17726 6566 17835 6568
rect 17769 6563 17835 6566
rect 4699 6560 5015 6561
rect 4699 6496 4705 6560
rect 4769 6496 4785 6560
rect 4849 6496 4865 6560
rect 4929 6496 4945 6560
rect 5009 6496 5015 6560
rect 4699 6495 5015 6496
rect 10886 6560 11202 6561
rect 10886 6496 10892 6560
rect 10956 6496 10972 6560
rect 11036 6496 11052 6560
rect 11116 6496 11132 6560
rect 11196 6496 11202 6560
rect 10886 6495 11202 6496
rect 17073 6560 17389 6561
rect 17073 6496 17079 6560
rect 17143 6496 17159 6560
rect 17223 6496 17239 6560
rect 17303 6496 17319 6560
rect 17383 6496 17389 6560
rect 17073 6495 17389 6496
rect 23260 6560 23576 6561
rect 23260 6496 23266 6560
rect 23330 6496 23346 6560
rect 23410 6496 23426 6560
rect 23490 6496 23506 6560
rect 23570 6496 23576 6560
rect 23260 6495 23576 6496
rect 9673 6354 9739 6357
rect 15745 6354 15811 6357
rect 17953 6354 18019 6357
rect 9673 6352 18019 6354
rect 9673 6296 9678 6352
rect 9734 6296 15750 6352
rect 15806 6296 17958 6352
rect 18014 6296 18019 6352
rect 9673 6294 18019 6296
rect 9673 6291 9739 6294
rect 15745 6291 15811 6294
rect 17953 6291 18019 6294
rect 5717 6218 5783 6221
rect 7925 6218 7991 6221
rect 9581 6218 9647 6221
rect 5717 6216 9647 6218
rect 5717 6160 5722 6216
rect 5778 6160 7930 6216
rect 7986 6160 9586 6216
rect 9642 6160 9647 6216
rect 5717 6158 9647 6160
rect 5717 6155 5783 6158
rect 7925 6155 7991 6158
rect 9581 6155 9647 6158
rect 25405 6218 25471 6221
rect 26237 6218 27037 6248
rect 25405 6216 27037 6218
rect 25405 6160 25410 6216
rect 25466 6160 27037 6216
rect 25405 6158 27037 6160
rect 25405 6155 25471 6158
rect 26237 6128 27037 6158
rect 4039 6016 4355 6017
rect 4039 5952 4045 6016
rect 4109 5952 4125 6016
rect 4189 5952 4205 6016
rect 4269 5952 4285 6016
rect 4349 5952 4355 6016
rect 4039 5951 4355 5952
rect 10226 6016 10542 6017
rect 10226 5952 10232 6016
rect 10296 5952 10312 6016
rect 10376 5952 10392 6016
rect 10456 5952 10472 6016
rect 10536 5952 10542 6016
rect 10226 5951 10542 5952
rect 16413 6016 16729 6017
rect 16413 5952 16419 6016
rect 16483 5952 16499 6016
rect 16563 5952 16579 6016
rect 16643 5952 16659 6016
rect 16723 5952 16729 6016
rect 16413 5951 16729 5952
rect 22600 6016 22916 6017
rect 22600 5952 22606 6016
rect 22670 5952 22686 6016
rect 22750 5952 22766 6016
rect 22830 5952 22846 6016
rect 22910 5952 22916 6016
rect 22600 5951 22916 5952
rect 16297 5674 16363 5677
rect 17125 5674 17191 5677
rect 16297 5672 17191 5674
rect 16297 5616 16302 5672
rect 16358 5616 17130 5672
rect 17186 5616 17191 5672
rect 16297 5614 17191 5616
rect 16297 5611 16363 5614
rect 17125 5611 17191 5614
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 4699 5472 5015 5473
rect 4699 5408 4705 5472
rect 4769 5408 4785 5472
rect 4849 5408 4865 5472
rect 4929 5408 4945 5472
rect 5009 5408 5015 5472
rect 4699 5407 5015 5408
rect 10886 5472 11202 5473
rect 10886 5408 10892 5472
rect 10956 5408 10972 5472
rect 11036 5408 11052 5472
rect 11116 5408 11132 5472
rect 11196 5408 11202 5472
rect 10886 5407 11202 5408
rect 17073 5472 17389 5473
rect 17073 5408 17079 5472
rect 17143 5408 17159 5472
rect 17223 5408 17239 5472
rect 17303 5408 17319 5472
rect 17383 5408 17389 5472
rect 17073 5407 17389 5408
rect 23260 5472 23576 5473
rect 23260 5408 23266 5472
rect 23330 5408 23346 5472
rect 23410 5408 23426 5472
rect 23490 5408 23506 5472
rect 23570 5408 23576 5472
rect 23260 5407 23576 5408
rect 14457 5266 14523 5269
rect 16021 5266 16087 5269
rect 14457 5264 16087 5266
rect 14457 5208 14462 5264
rect 14518 5208 16026 5264
rect 16082 5208 16087 5264
rect 14457 5206 16087 5208
rect 14457 5203 14523 5206
rect 16021 5203 16087 5206
rect 4039 4928 4355 4929
rect 0 4858 800 4888
rect 4039 4864 4045 4928
rect 4109 4864 4125 4928
rect 4189 4864 4205 4928
rect 4269 4864 4285 4928
rect 4349 4864 4355 4928
rect 4039 4863 4355 4864
rect 10226 4928 10542 4929
rect 10226 4864 10232 4928
rect 10296 4864 10312 4928
rect 10376 4864 10392 4928
rect 10456 4864 10472 4928
rect 10536 4864 10542 4928
rect 10226 4863 10542 4864
rect 16413 4928 16729 4929
rect 16413 4864 16419 4928
rect 16483 4864 16499 4928
rect 16563 4864 16579 4928
rect 16643 4864 16659 4928
rect 16723 4864 16729 4928
rect 16413 4863 16729 4864
rect 22600 4928 22916 4929
rect 22600 4864 22606 4928
rect 22670 4864 22686 4928
rect 22750 4864 22766 4928
rect 22830 4864 22846 4928
rect 22910 4864 22916 4928
rect 22600 4863 22916 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 25405 4858 25471 4861
rect 26237 4858 27037 4888
rect 25405 4856 27037 4858
rect 25405 4800 25410 4856
rect 25466 4800 27037 4856
rect 25405 4798 27037 4800
rect 25405 4795 25471 4798
rect 26237 4768 27037 4798
rect 15561 4722 15627 4725
rect 16389 4722 16455 4725
rect 15561 4720 16455 4722
rect 15561 4664 15566 4720
rect 15622 4664 16394 4720
rect 16450 4664 16455 4720
rect 15561 4662 16455 4664
rect 15561 4659 15627 4662
rect 16389 4659 16455 4662
rect 1577 4586 1643 4589
rect 21081 4586 21147 4589
rect 1577 4584 21147 4586
rect 1577 4528 1582 4584
rect 1638 4528 21086 4584
rect 21142 4528 21147 4584
rect 1577 4526 21147 4528
rect 1577 4523 1643 4526
rect 21081 4523 21147 4526
rect 4699 4384 5015 4385
rect 4699 4320 4705 4384
rect 4769 4320 4785 4384
rect 4849 4320 4865 4384
rect 4929 4320 4945 4384
rect 5009 4320 5015 4384
rect 4699 4319 5015 4320
rect 10886 4384 11202 4385
rect 10886 4320 10892 4384
rect 10956 4320 10972 4384
rect 11036 4320 11052 4384
rect 11116 4320 11132 4384
rect 11196 4320 11202 4384
rect 10886 4319 11202 4320
rect 17073 4384 17389 4385
rect 17073 4320 17079 4384
rect 17143 4320 17159 4384
rect 17223 4320 17239 4384
rect 17303 4320 17319 4384
rect 17383 4320 17389 4384
rect 17073 4319 17389 4320
rect 23260 4384 23576 4385
rect 23260 4320 23266 4384
rect 23330 4320 23346 4384
rect 23410 4320 23426 4384
rect 23490 4320 23506 4384
rect 23570 4320 23576 4384
rect 23260 4319 23576 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 25405 4178 25471 4181
rect 26237 4178 27037 4208
rect 25405 4176 27037 4178
rect 25405 4120 25410 4176
rect 25466 4120 27037 4176
rect 25405 4118 27037 4120
rect 25405 4115 25471 4118
rect 26237 4088 27037 4118
rect 4039 3840 4355 3841
rect 4039 3776 4045 3840
rect 4109 3776 4125 3840
rect 4189 3776 4205 3840
rect 4269 3776 4285 3840
rect 4349 3776 4355 3840
rect 4039 3775 4355 3776
rect 10226 3840 10542 3841
rect 10226 3776 10232 3840
rect 10296 3776 10312 3840
rect 10376 3776 10392 3840
rect 10456 3776 10472 3840
rect 10536 3776 10542 3840
rect 10226 3775 10542 3776
rect 16413 3840 16729 3841
rect 16413 3776 16419 3840
rect 16483 3776 16499 3840
rect 16563 3776 16579 3840
rect 16643 3776 16659 3840
rect 16723 3776 16729 3840
rect 16413 3775 16729 3776
rect 22600 3840 22916 3841
rect 22600 3776 22606 3840
rect 22670 3776 22686 3840
rect 22750 3776 22766 3840
rect 22830 3776 22846 3840
rect 22910 3776 22916 3840
rect 22600 3775 22916 3776
rect 0 3498 800 3528
rect 1025 3498 1091 3501
rect 0 3496 1091 3498
rect 0 3440 1030 3496
rect 1086 3440 1091 3496
rect 0 3438 1091 3440
rect 0 3408 800 3438
rect 1025 3435 1091 3438
rect 25957 3498 26023 3501
rect 26237 3498 27037 3528
rect 25957 3496 27037 3498
rect 25957 3440 25962 3496
rect 26018 3440 27037 3496
rect 25957 3438 27037 3440
rect 25957 3435 26023 3438
rect 26237 3408 27037 3438
rect 4699 3296 5015 3297
rect 4699 3232 4705 3296
rect 4769 3232 4785 3296
rect 4849 3232 4865 3296
rect 4929 3232 4945 3296
rect 5009 3232 5015 3296
rect 4699 3231 5015 3232
rect 10886 3296 11202 3297
rect 10886 3232 10892 3296
rect 10956 3232 10972 3296
rect 11036 3232 11052 3296
rect 11116 3232 11132 3296
rect 11196 3232 11202 3296
rect 10886 3231 11202 3232
rect 17073 3296 17389 3297
rect 17073 3232 17079 3296
rect 17143 3232 17159 3296
rect 17223 3232 17239 3296
rect 17303 3232 17319 3296
rect 17383 3232 17389 3296
rect 17073 3231 17389 3232
rect 23260 3296 23576 3297
rect 23260 3232 23266 3296
rect 23330 3232 23346 3296
rect 23410 3232 23426 3296
rect 23490 3232 23506 3296
rect 23570 3232 23576 3296
rect 23260 3231 23576 3232
rect 2037 3090 2103 3093
rect 21081 3090 21147 3093
rect 2037 3088 21147 3090
rect 2037 3032 2042 3088
rect 2098 3032 21086 3088
rect 21142 3032 21147 3088
rect 2037 3030 21147 3032
rect 2037 3027 2103 3030
rect 21081 3027 21147 3030
rect 9857 2954 9923 2957
rect 12801 2954 12867 2957
rect 9857 2952 12867 2954
rect 9857 2896 9862 2952
rect 9918 2896 12806 2952
rect 12862 2896 12867 2952
rect 9857 2894 12867 2896
rect 9857 2891 9923 2894
rect 12801 2891 12867 2894
rect 25129 2818 25195 2821
rect 26237 2818 27037 2848
rect 25129 2816 27037 2818
rect 25129 2760 25134 2816
rect 25190 2760 27037 2816
rect 25129 2758 27037 2760
rect 25129 2755 25195 2758
rect 4039 2752 4355 2753
rect 4039 2688 4045 2752
rect 4109 2688 4125 2752
rect 4189 2688 4205 2752
rect 4269 2688 4285 2752
rect 4349 2688 4355 2752
rect 4039 2687 4355 2688
rect 10226 2752 10542 2753
rect 10226 2688 10232 2752
rect 10296 2688 10312 2752
rect 10376 2688 10392 2752
rect 10456 2688 10472 2752
rect 10536 2688 10542 2752
rect 10226 2687 10542 2688
rect 16413 2752 16729 2753
rect 16413 2688 16419 2752
rect 16483 2688 16499 2752
rect 16563 2688 16579 2752
rect 16643 2688 16659 2752
rect 16723 2688 16729 2752
rect 16413 2687 16729 2688
rect 22600 2752 22916 2753
rect 22600 2688 22606 2752
rect 22670 2688 22686 2752
rect 22750 2688 22766 2752
rect 22830 2688 22846 2752
rect 22910 2688 22916 2752
rect 26237 2728 27037 2758
rect 22600 2687 22916 2688
rect 15193 2682 15259 2685
rect 15326 2682 15332 2684
rect 15193 2680 15332 2682
rect 15193 2624 15198 2680
rect 15254 2624 15332 2680
rect 15193 2622 15332 2624
rect 15193 2619 15259 2622
rect 15326 2620 15332 2622
rect 15396 2620 15402 2684
rect 3877 2410 3943 2413
rect 19425 2410 19491 2413
rect 3877 2408 19491 2410
rect 3877 2352 3882 2408
rect 3938 2352 19430 2408
rect 19486 2352 19491 2408
rect 3877 2350 19491 2352
rect 3877 2347 3943 2350
rect 19425 2347 19491 2350
rect 4699 2208 5015 2209
rect 0 2138 800 2168
rect 4699 2144 4705 2208
rect 4769 2144 4785 2208
rect 4849 2144 4865 2208
rect 4929 2144 4945 2208
rect 5009 2144 5015 2208
rect 4699 2143 5015 2144
rect 10886 2208 11202 2209
rect 10886 2144 10892 2208
rect 10956 2144 10972 2208
rect 11036 2144 11052 2208
rect 11116 2144 11132 2208
rect 11196 2144 11202 2208
rect 10886 2143 11202 2144
rect 17073 2208 17389 2209
rect 17073 2144 17079 2208
rect 17143 2144 17159 2208
rect 17223 2144 17239 2208
rect 17303 2144 17319 2208
rect 17383 2144 17389 2208
rect 17073 2143 17389 2144
rect 23260 2208 23576 2209
rect 23260 2144 23266 2208
rect 23330 2144 23346 2208
rect 23410 2144 23426 2208
rect 23490 2144 23506 2208
rect 23570 2144 23576 2208
rect 23260 2143 23576 2144
rect 1577 2138 1643 2141
rect 0 2136 1643 2138
rect 0 2080 1582 2136
rect 1638 2080 1643 2136
rect 0 2078 1643 2080
rect 0 2048 800 2078
rect 1577 2075 1643 2078
rect 0 1458 800 1488
rect 1301 1458 1367 1461
rect 0 1456 1367 1458
rect 0 1400 1306 1456
rect 1362 1400 1367 1456
rect 0 1398 1367 1400
rect 0 1368 800 1398
rect 1301 1395 1367 1398
rect 24669 1458 24735 1461
rect 26237 1458 27037 1488
rect 24669 1456 27037 1458
rect 24669 1400 24674 1456
rect 24730 1400 27037 1456
rect 24669 1398 27037 1400
rect 24669 1395 24735 1398
rect 26237 1368 27037 1398
rect 25037 914 25103 917
rect 25037 912 25146 914
rect 25037 856 25042 912
rect 25098 856 25146 912
rect 25037 851 25146 856
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 25086 778 25146 851
rect 26237 778 27037 808
rect 25086 718 27037 778
rect 0 688 800 718
rect 2773 715 2839 718
rect 26237 688 27037 718
rect 25865 98 25931 101
rect 26237 98 27037 128
rect 25865 96 27037 98
rect 25865 40 25870 96
rect 25926 40 27037 96
rect 25865 38 27037 40
rect 25865 35 25931 38
rect 26237 8 27037 38
<< via3 >>
rect 4045 26684 4109 26688
rect 4045 26628 4049 26684
rect 4049 26628 4105 26684
rect 4105 26628 4109 26684
rect 4045 26624 4109 26628
rect 4125 26684 4189 26688
rect 4125 26628 4129 26684
rect 4129 26628 4185 26684
rect 4185 26628 4189 26684
rect 4125 26624 4189 26628
rect 4205 26684 4269 26688
rect 4205 26628 4209 26684
rect 4209 26628 4265 26684
rect 4265 26628 4269 26684
rect 4205 26624 4269 26628
rect 4285 26684 4349 26688
rect 4285 26628 4289 26684
rect 4289 26628 4345 26684
rect 4345 26628 4349 26684
rect 4285 26624 4349 26628
rect 10232 26684 10296 26688
rect 10232 26628 10236 26684
rect 10236 26628 10292 26684
rect 10292 26628 10296 26684
rect 10232 26624 10296 26628
rect 10312 26684 10376 26688
rect 10312 26628 10316 26684
rect 10316 26628 10372 26684
rect 10372 26628 10376 26684
rect 10312 26624 10376 26628
rect 10392 26684 10456 26688
rect 10392 26628 10396 26684
rect 10396 26628 10452 26684
rect 10452 26628 10456 26684
rect 10392 26624 10456 26628
rect 10472 26684 10536 26688
rect 10472 26628 10476 26684
rect 10476 26628 10532 26684
rect 10532 26628 10536 26684
rect 10472 26624 10536 26628
rect 16419 26684 16483 26688
rect 16419 26628 16423 26684
rect 16423 26628 16479 26684
rect 16479 26628 16483 26684
rect 16419 26624 16483 26628
rect 16499 26684 16563 26688
rect 16499 26628 16503 26684
rect 16503 26628 16559 26684
rect 16559 26628 16563 26684
rect 16499 26624 16563 26628
rect 16579 26684 16643 26688
rect 16579 26628 16583 26684
rect 16583 26628 16639 26684
rect 16639 26628 16643 26684
rect 16579 26624 16643 26628
rect 16659 26684 16723 26688
rect 16659 26628 16663 26684
rect 16663 26628 16719 26684
rect 16719 26628 16723 26684
rect 16659 26624 16723 26628
rect 22606 26684 22670 26688
rect 22606 26628 22610 26684
rect 22610 26628 22666 26684
rect 22666 26628 22670 26684
rect 22606 26624 22670 26628
rect 22686 26684 22750 26688
rect 22686 26628 22690 26684
rect 22690 26628 22746 26684
rect 22746 26628 22750 26684
rect 22686 26624 22750 26628
rect 22766 26684 22830 26688
rect 22766 26628 22770 26684
rect 22770 26628 22826 26684
rect 22826 26628 22830 26684
rect 22766 26624 22830 26628
rect 22846 26684 22910 26688
rect 22846 26628 22850 26684
rect 22850 26628 22906 26684
rect 22906 26628 22910 26684
rect 22846 26624 22910 26628
rect 4705 26140 4769 26144
rect 4705 26084 4709 26140
rect 4709 26084 4765 26140
rect 4765 26084 4769 26140
rect 4705 26080 4769 26084
rect 4785 26140 4849 26144
rect 4785 26084 4789 26140
rect 4789 26084 4845 26140
rect 4845 26084 4849 26140
rect 4785 26080 4849 26084
rect 4865 26140 4929 26144
rect 4865 26084 4869 26140
rect 4869 26084 4925 26140
rect 4925 26084 4929 26140
rect 4865 26080 4929 26084
rect 4945 26140 5009 26144
rect 4945 26084 4949 26140
rect 4949 26084 5005 26140
rect 5005 26084 5009 26140
rect 4945 26080 5009 26084
rect 10892 26140 10956 26144
rect 10892 26084 10896 26140
rect 10896 26084 10952 26140
rect 10952 26084 10956 26140
rect 10892 26080 10956 26084
rect 10972 26140 11036 26144
rect 10972 26084 10976 26140
rect 10976 26084 11032 26140
rect 11032 26084 11036 26140
rect 10972 26080 11036 26084
rect 11052 26140 11116 26144
rect 11052 26084 11056 26140
rect 11056 26084 11112 26140
rect 11112 26084 11116 26140
rect 11052 26080 11116 26084
rect 11132 26140 11196 26144
rect 11132 26084 11136 26140
rect 11136 26084 11192 26140
rect 11192 26084 11196 26140
rect 11132 26080 11196 26084
rect 17079 26140 17143 26144
rect 17079 26084 17083 26140
rect 17083 26084 17139 26140
rect 17139 26084 17143 26140
rect 17079 26080 17143 26084
rect 17159 26140 17223 26144
rect 17159 26084 17163 26140
rect 17163 26084 17219 26140
rect 17219 26084 17223 26140
rect 17159 26080 17223 26084
rect 17239 26140 17303 26144
rect 17239 26084 17243 26140
rect 17243 26084 17299 26140
rect 17299 26084 17303 26140
rect 17239 26080 17303 26084
rect 17319 26140 17383 26144
rect 17319 26084 17323 26140
rect 17323 26084 17379 26140
rect 17379 26084 17383 26140
rect 17319 26080 17383 26084
rect 23266 26140 23330 26144
rect 23266 26084 23270 26140
rect 23270 26084 23326 26140
rect 23326 26084 23330 26140
rect 23266 26080 23330 26084
rect 23346 26140 23410 26144
rect 23346 26084 23350 26140
rect 23350 26084 23406 26140
rect 23406 26084 23410 26140
rect 23346 26080 23410 26084
rect 23426 26140 23490 26144
rect 23426 26084 23430 26140
rect 23430 26084 23486 26140
rect 23486 26084 23490 26140
rect 23426 26080 23490 26084
rect 23506 26140 23570 26144
rect 23506 26084 23510 26140
rect 23510 26084 23566 26140
rect 23566 26084 23570 26140
rect 23506 26080 23570 26084
rect 4045 25596 4109 25600
rect 4045 25540 4049 25596
rect 4049 25540 4105 25596
rect 4105 25540 4109 25596
rect 4045 25536 4109 25540
rect 4125 25596 4189 25600
rect 4125 25540 4129 25596
rect 4129 25540 4185 25596
rect 4185 25540 4189 25596
rect 4125 25536 4189 25540
rect 4205 25596 4269 25600
rect 4205 25540 4209 25596
rect 4209 25540 4265 25596
rect 4265 25540 4269 25596
rect 4205 25536 4269 25540
rect 4285 25596 4349 25600
rect 4285 25540 4289 25596
rect 4289 25540 4345 25596
rect 4345 25540 4349 25596
rect 4285 25536 4349 25540
rect 10232 25596 10296 25600
rect 10232 25540 10236 25596
rect 10236 25540 10292 25596
rect 10292 25540 10296 25596
rect 10232 25536 10296 25540
rect 10312 25596 10376 25600
rect 10312 25540 10316 25596
rect 10316 25540 10372 25596
rect 10372 25540 10376 25596
rect 10312 25536 10376 25540
rect 10392 25596 10456 25600
rect 10392 25540 10396 25596
rect 10396 25540 10452 25596
rect 10452 25540 10456 25596
rect 10392 25536 10456 25540
rect 10472 25596 10536 25600
rect 10472 25540 10476 25596
rect 10476 25540 10532 25596
rect 10532 25540 10536 25596
rect 10472 25536 10536 25540
rect 16419 25596 16483 25600
rect 16419 25540 16423 25596
rect 16423 25540 16479 25596
rect 16479 25540 16483 25596
rect 16419 25536 16483 25540
rect 16499 25596 16563 25600
rect 16499 25540 16503 25596
rect 16503 25540 16559 25596
rect 16559 25540 16563 25596
rect 16499 25536 16563 25540
rect 16579 25596 16643 25600
rect 16579 25540 16583 25596
rect 16583 25540 16639 25596
rect 16639 25540 16643 25596
rect 16579 25536 16643 25540
rect 16659 25596 16723 25600
rect 16659 25540 16663 25596
rect 16663 25540 16719 25596
rect 16719 25540 16723 25596
rect 16659 25536 16723 25540
rect 22606 25596 22670 25600
rect 22606 25540 22610 25596
rect 22610 25540 22666 25596
rect 22666 25540 22670 25596
rect 22606 25536 22670 25540
rect 22686 25596 22750 25600
rect 22686 25540 22690 25596
rect 22690 25540 22746 25596
rect 22746 25540 22750 25596
rect 22686 25536 22750 25540
rect 22766 25596 22830 25600
rect 22766 25540 22770 25596
rect 22770 25540 22826 25596
rect 22826 25540 22830 25596
rect 22766 25536 22830 25540
rect 22846 25596 22910 25600
rect 22846 25540 22850 25596
rect 22850 25540 22906 25596
rect 22906 25540 22910 25596
rect 22846 25536 22910 25540
rect 4705 25052 4769 25056
rect 4705 24996 4709 25052
rect 4709 24996 4765 25052
rect 4765 24996 4769 25052
rect 4705 24992 4769 24996
rect 4785 25052 4849 25056
rect 4785 24996 4789 25052
rect 4789 24996 4845 25052
rect 4845 24996 4849 25052
rect 4785 24992 4849 24996
rect 4865 25052 4929 25056
rect 4865 24996 4869 25052
rect 4869 24996 4925 25052
rect 4925 24996 4929 25052
rect 4865 24992 4929 24996
rect 4945 25052 5009 25056
rect 4945 24996 4949 25052
rect 4949 24996 5005 25052
rect 5005 24996 5009 25052
rect 4945 24992 5009 24996
rect 10892 25052 10956 25056
rect 10892 24996 10896 25052
rect 10896 24996 10952 25052
rect 10952 24996 10956 25052
rect 10892 24992 10956 24996
rect 10972 25052 11036 25056
rect 10972 24996 10976 25052
rect 10976 24996 11032 25052
rect 11032 24996 11036 25052
rect 10972 24992 11036 24996
rect 11052 25052 11116 25056
rect 11052 24996 11056 25052
rect 11056 24996 11112 25052
rect 11112 24996 11116 25052
rect 11052 24992 11116 24996
rect 11132 25052 11196 25056
rect 11132 24996 11136 25052
rect 11136 24996 11192 25052
rect 11192 24996 11196 25052
rect 11132 24992 11196 24996
rect 17079 25052 17143 25056
rect 17079 24996 17083 25052
rect 17083 24996 17139 25052
rect 17139 24996 17143 25052
rect 17079 24992 17143 24996
rect 17159 25052 17223 25056
rect 17159 24996 17163 25052
rect 17163 24996 17219 25052
rect 17219 24996 17223 25052
rect 17159 24992 17223 24996
rect 17239 25052 17303 25056
rect 17239 24996 17243 25052
rect 17243 24996 17299 25052
rect 17299 24996 17303 25052
rect 17239 24992 17303 24996
rect 17319 25052 17383 25056
rect 17319 24996 17323 25052
rect 17323 24996 17379 25052
rect 17379 24996 17383 25052
rect 17319 24992 17383 24996
rect 23266 25052 23330 25056
rect 23266 24996 23270 25052
rect 23270 24996 23326 25052
rect 23326 24996 23330 25052
rect 23266 24992 23330 24996
rect 23346 25052 23410 25056
rect 23346 24996 23350 25052
rect 23350 24996 23406 25052
rect 23406 24996 23410 25052
rect 23346 24992 23410 24996
rect 23426 25052 23490 25056
rect 23426 24996 23430 25052
rect 23430 24996 23486 25052
rect 23486 24996 23490 25052
rect 23426 24992 23490 24996
rect 23506 25052 23570 25056
rect 23506 24996 23510 25052
rect 23510 24996 23566 25052
rect 23566 24996 23570 25052
rect 23506 24992 23570 24996
rect 9812 24652 9876 24716
rect 4045 24508 4109 24512
rect 4045 24452 4049 24508
rect 4049 24452 4105 24508
rect 4105 24452 4109 24508
rect 4045 24448 4109 24452
rect 4125 24508 4189 24512
rect 4125 24452 4129 24508
rect 4129 24452 4185 24508
rect 4185 24452 4189 24508
rect 4125 24448 4189 24452
rect 4205 24508 4269 24512
rect 4205 24452 4209 24508
rect 4209 24452 4265 24508
rect 4265 24452 4269 24508
rect 4205 24448 4269 24452
rect 4285 24508 4349 24512
rect 4285 24452 4289 24508
rect 4289 24452 4345 24508
rect 4345 24452 4349 24508
rect 4285 24448 4349 24452
rect 10232 24508 10296 24512
rect 10232 24452 10236 24508
rect 10236 24452 10292 24508
rect 10292 24452 10296 24508
rect 10232 24448 10296 24452
rect 10312 24508 10376 24512
rect 10312 24452 10316 24508
rect 10316 24452 10372 24508
rect 10372 24452 10376 24508
rect 10312 24448 10376 24452
rect 10392 24508 10456 24512
rect 10392 24452 10396 24508
rect 10396 24452 10452 24508
rect 10452 24452 10456 24508
rect 10392 24448 10456 24452
rect 10472 24508 10536 24512
rect 10472 24452 10476 24508
rect 10476 24452 10532 24508
rect 10532 24452 10536 24508
rect 10472 24448 10536 24452
rect 16419 24508 16483 24512
rect 16419 24452 16423 24508
rect 16423 24452 16479 24508
rect 16479 24452 16483 24508
rect 16419 24448 16483 24452
rect 16499 24508 16563 24512
rect 16499 24452 16503 24508
rect 16503 24452 16559 24508
rect 16559 24452 16563 24508
rect 16499 24448 16563 24452
rect 16579 24508 16643 24512
rect 16579 24452 16583 24508
rect 16583 24452 16639 24508
rect 16639 24452 16643 24508
rect 16579 24448 16643 24452
rect 16659 24508 16723 24512
rect 16659 24452 16663 24508
rect 16663 24452 16719 24508
rect 16719 24452 16723 24508
rect 16659 24448 16723 24452
rect 22606 24508 22670 24512
rect 22606 24452 22610 24508
rect 22610 24452 22666 24508
rect 22666 24452 22670 24508
rect 22606 24448 22670 24452
rect 22686 24508 22750 24512
rect 22686 24452 22690 24508
rect 22690 24452 22746 24508
rect 22746 24452 22750 24508
rect 22686 24448 22750 24452
rect 22766 24508 22830 24512
rect 22766 24452 22770 24508
rect 22770 24452 22826 24508
rect 22826 24452 22830 24508
rect 22766 24448 22830 24452
rect 22846 24508 22910 24512
rect 22846 24452 22850 24508
rect 22850 24452 22906 24508
rect 22906 24452 22910 24508
rect 22846 24448 22910 24452
rect 4705 23964 4769 23968
rect 4705 23908 4709 23964
rect 4709 23908 4765 23964
rect 4765 23908 4769 23964
rect 4705 23904 4769 23908
rect 4785 23964 4849 23968
rect 4785 23908 4789 23964
rect 4789 23908 4845 23964
rect 4845 23908 4849 23964
rect 4785 23904 4849 23908
rect 4865 23964 4929 23968
rect 4865 23908 4869 23964
rect 4869 23908 4925 23964
rect 4925 23908 4929 23964
rect 4865 23904 4929 23908
rect 4945 23964 5009 23968
rect 4945 23908 4949 23964
rect 4949 23908 5005 23964
rect 5005 23908 5009 23964
rect 4945 23904 5009 23908
rect 10892 23964 10956 23968
rect 10892 23908 10896 23964
rect 10896 23908 10952 23964
rect 10952 23908 10956 23964
rect 10892 23904 10956 23908
rect 10972 23964 11036 23968
rect 10972 23908 10976 23964
rect 10976 23908 11032 23964
rect 11032 23908 11036 23964
rect 10972 23904 11036 23908
rect 11052 23964 11116 23968
rect 11052 23908 11056 23964
rect 11056 23908 11112 23964
rect 11112 23908 11116 23964
rect 11052 23904 11116 23908
rect 11132 23964 11196 23968
rect 11132 23908 11136 23964
rect 11136 23908 11192 23964
rect 11192 23908 11196 23964
rect 11132 23904 11196 23908
rect 17079 23964 17143 23968
rect 17079 23908 17083 23964
rect 17083 23908 17139 23964
rect 17139 23908 17143 23964
rect 17079 23904 17143 23908
rect 17159 23964 17223 23968
rect 17159 23908 17163 23964
rect 17163 23908 17219 23964
rect 17219 23908 17223 23964
rect 17159 23904 17223 23908
rect 17239 23964 17303 23968
rect 17239 23908 17243 23964
rect 17243 23908 17299 23964
rect 17299 23908 17303 23964
rect 17239 23904 17303 23908
rect 17319 23964 17383 23968
rect 17319 23908 17323 23964
rect 17323 23908 17379 23964
rect 17379 23908 17383 23964
rect 17319 23904 17383 23908
rect 23266 23964 23330 23968
rect 23266 23908 23270 23964
rect 23270 23908 23326 23964
rect 23326 23908 23330 23964
rect 23266 23904 23330 23908
rect 23346 23964 23410 23968
rect 23346 23908 23350 23964
rect 23350 23908 23406 23964
rect 23406 23908 23410 23964
rect 23346 23904 23410 23908
rect 23426 23964 23490 23968
rect 23426 23908 23430 23964
rect 23430 23908 23486 23964
rect 23486 23908 23490 23964
rect 23426 23904 23490 23908
rect 23506 23964 23570 23968
rect 23506 23908 23510 23964
rect 23510 23908 23566 23964
rect 23566 23908 23570 23964
rect 23506 23904 23570 23908
rect 4045 23420 4109 23424
rect 4045 23364 4049 23420
rect 4049 23364 4105 23420
rect 4105 23364 4109 23420
rect 4045 23360 4109 23364
rect 4125 23420 4189 23424
rect 4125 23364 4129 23420
rect 4129 23364 4185 23420
rect 4185 23364 4189 23420
rect 4125 23360 4189 23364
rect 4205 23420 4269 23424
rect 4205 23364 4209 23420
rect 4209 23364 4265 23420
rect 4265 23364 4269 23420
rect 4205 23360 4269 23364
rect 4285 23420 4349 23424
rect 4285 23364 4289 23420
rect 4289 23364 4345 23420
rect 4345 23364 4349 23420
rect 4285 23360 4349 23364
rect 10232 23420 10296 23424
rect 10232 23364 10236 23420
rect 10236 23364 10292 23420
rect 10292 23364 10296 23420
rect 10232 23360 10296 23364
rect 10312 23420 10376 23424
rect 10312 23364 10316 23420
rect 10316 23364 10372 23420
rect 10372 23364 10376 23420
rect 10312 23360 10376 23364
rect 10392 23420 10456 23424
rect 10392 23364 10396 23420
rect 10396 23364 10452 23420
rect 10452 23364 10456 23420
rect 10392 23360 10456 23364
rect 10472 23420 10536 23424
rect 10472 23364 10476 23420
rect 10476 23364 10532 23420
rect 10532 23364 10536 23420
rect 10472 23360 10536 23364
rect 16419 23420 16483 23424
rect 16419 23364 16423 23420
rect 16423 23364 16479 23420
rect 16479 23364 16483 23420
rect 16419 23360 16483 23364
rect 16499 23420 16563 23424
rect 16499 23364 16503 23420
rect 16503 23364 16559 23420
rect 16559 23364 16563 23420
rect 16499 23360 16563 23364
rect 16579 23420 16643 23424
rect 16579 23364 16583 23420
rect 16583 23364 16639 23420
rect 16639 23364 16643 23420
rect 16579 23360 16643 23364
rect 16659 23420 16723 23424
rect 16659 23364 16663 23420
rect 16663 23364 16719 23420
rect 16719 23364 16723 23420
rect 16659 23360 16723 23364
rect 22606 23420 22670 23424
rect 22606 23364 22610 23420
rect 22610 23364 22666 23420
rect 22666 23364 22670 23420
rect 22606 23360 22670 23364
rect 22686 23420 22750 23424
rect 22686 23364 22690 23420
rect 22690 23364 22746 23420
rect 22746 23364 22750 23420
rect 22686 23360 22750 23364
rect 22766 23420 22830 23424
rect 22766 23364 22770 23420
rect 22770 23364 22826 23420
rect 22826 23364 22830 23420
rect 22766 23360 22830 23364
rect 22846 23420 22910 23424
rect 22846 23364 22850 23420
rect 22850 23364 22906 23420
rect 22906 23364 22910 23420
rect 22846 23360 22910 23364
rect 4705 22876 4769 22880
rect 4705 22820 4709 22876
rect 4709 22820 4765 22876
rect 4765 22820 4769 22876
rect 4705 22816 4769 22820
rect 4785 22876 4849 22880
rect 4785 22820 4789 22876
rect 4789 22820 4845 22876
rect 4845 22820 4849 22876
rect 4785 22816 4849 22820
rect 4865 22876 4929 22880
rect 4865 22820 4869 22876
rect 4869 22820 4925 22876
rect 4925 22820 4929 22876
rect 4865 22816 4929 22820
rect 4945 22876 5009 22880
rect 4945 22820 4949 22876
rect 4949 22820 5005 22876
rect 5005 22820 5009 22876
rect 4945 22816 5009 22820
rect 10892 22876 10956 22880
rect 10892 22820 10896 22876
rect 10896 22820 10952 22876
rect 10952 22820 10956 22876
rect 10892 22816 10956 22820
rect 10972 22876 11036 22880
rect 10972 22820 10976 22876
rect 10976 22820 11032 22876
rect 11032 22820 11036 22876
rect 10972 22816 11036 22820
rect 11052 22876 11116 22880
rect 11052 22820 11056 22876
rect 11056 22820 11112 22876
rect 11112 22820 11116 22876
rect 11052 22816 11116 22820
rect 11132 22876 11196 22880
rect 11132 22820 11136 22876
rect 11136 22820 11192 22876
rect 11192 22820 11196 22876
rect 11132 22816 11196 22820
rect 17079 22876 17143 22880
rect 17079 22820 17083 22876
rect 17083 22820 17139 22876
rect 17139 22820 17143 22876
rect 17079 22816 17143 22820
rect 17159 22876 17223 22880
rect 17159 22820 17163 22876
rect 17163 22820 17219 22876
rect 17219 22820 17223 22876
rect 17159 22816 17223 22820
rect 17239 22876 17303 22880
rect 17239 22820 17243 22876
rect 17243 22820 17299 22876
rect 17299 22820 17303 22876
rect 17239 22816 17303 22820
rect 17319 22876 17383 22880
rect 17319 22820 17323 22876
rect 17323 22820 17379 22876
rect 17379 22820 17383 22876
rect 17319 22816 17383 22820
rect 23266 22876 23330 22880
rect 23266 22820 23270 22876
rect 23270 22820 23326 22876
rect 23326 22820 23330 22876
rect 23266 22816 23330 22820
rect 23346 22876 23410 22880
rect 23346 22820 23350 22876
rect 23350 22820 23406 22876
rect 23406 22820 23410 22876
rect 23346 22816 23410 22820
rect 23426 22876 23490 22880
rect 23426 22820 23430 22876
rect 23430 22820 23486 22876
rect 23486 22820 23490 22876
rect 23426 22816 23490 22820
rect 23506 22876 23570 22880
rect 23506 22820 23510 22876
rect 23510 22820 23566 22876
rect 23566 22820 23570 22876
rect 23506 22816 23570 22820
rect 9812 22808 9876 22812
rect 9812 22752 9826 22808
rect 9826 22752 9876 22808
rect 9812 22748 9876 22752
rect 4045 22332 4109 22336
rect 4045 22276 4049 22332
rect 4049 22276 4105 22332
rect 4105 22276 4109 22332
rect 4045 22272 4109 22276
rect 4125 22332 4189 22336
rect 4125 22276 4129 22332
rect 4129 22276 4185 22332
rect 4185 22276 4189 22332
rect 4125 22272 4189 22276
rect 4205 22332 4269 22336
rect 4205 22276 4209 22332
rect 4209 22276 4265 22332
rect 4265 22276 4269 22332
rect 4205 22272 4269 22276
rect 4285 22332 4349 22336
rect 4285 22276 4289 22332
rect 4289 22276 4345 22332
rect 4345 22276 4349 22332
rect 4285 22272 4349 22276
rect 10232 22332 10296 22336
rect 10232 22276 10236 22332
rect 10236 22276 10292 22332
rect 10292 22276 10296 22332
rect 10232 22272 10296 22276
rect 10312 22332 10376 22336
rect 10312 22276 10316 22332
rect 10316 22276 10372 22332
rect 10372 22276 10376 22332
rect 10312 22272 10376 22276
rect 10392 22332 10456 22336
rect 10392 22276 10396 22332
rect 10396 22276 10452 22332
rect 10452 22276 10456 22332
rect 10392 22272 10456 22276
rect 10472 22332 10536 22336
rect 10472 22276 10476 22332
rect 10476 22276 10532 22332
rect 10532 22276 10536 22332
rect 10472 22272 10536 22276
rect 16419 22332 16483 22336
rect 16419 22276 16423 22332
rect 16423 22276 16479 22332
rect 16479 22276 16483 22332
rect 16419 22272 16483 22276
rect 16499 22332 16563 22336
rect 16499 22276 16503 22332
rect 16503 22276 16559 22332
rect 16559 22276 16563 22332
rect 16499 22272 16563 22276
rect 16579 22332 16643 22336
rect 16579 22276 16583 22332
rect 16583 22276 16639 22332
rect 16639 22276 16643 22332
rect 16579 22272 16643 22276
rect 16659 22332 16723 22336
rect 16659 22276 16663 22332
rect 16663 22276 16719 22332
rect 16719 22276 16723 22332
rect 16659 22272 16723 22276
rect 22606 22332 22670 22336
rect 22606 22276 22610 22332
rect 22610 22276 22666 22332
rect 22666 22276 22670 22332
rect 22606 22272 22670 22276
rect 22686 22332 22750 22336
rect 22686 22276 22690 22332
rect 22690 22276 22746 22332
rect 22746 22276 22750 22332
rect 22686 22272 22750 22276
rect 22766 22332 22830 22336
rect 22766 22276 22770 22332
rect 22770 22276 22826 22332
rect 22826 22276 22830 22332
rect 22766 22272 22830 22276
rect 22846 22332 22910 22336
rect 22846 22276 22850 22332
rect 22850 22276 22906 22332
rect 22906 22276 22910 22332
rect 22846 22272 22910 22276
rect 4705 21788 4769 21792
rect 4705 21732 4709 21788
rect 4709 21732 4765 21788
rect 4765 21732 4769 21788
rect 4705 21728 4769 21732
rect 4785 21788 4849 21792
rect 4785 21732 4789 21788
rect 4789 21732 4845 21788
rect 4845 21732 4849 21788
rect 4785 21728 4849 21732
rect 4865 21788 4929 21792
rect 4865 21732 4869 21788
rect 4869 21732 4925 21788
rect 4925 21732 4929 21788
rect 4865 21728 4929 21732
rect 4945 21788 5009 21792
rect 4945 21732 4949 21788
rect 4949 21732 5005 21788
rect 5005 21732 5009 21788
rect 4945 21728 5009 21732
rect 10892 21788 10956 21792
rect 10892 21732 10896 21788
rect 10896 21732 10952 21788
rect 10952 21732 10956 21788
rect 10892 21728 10956 21732
rect 10972 21788 11036 21792
rect 10972 21732 10976 21788
rect 10976 21732 11032 21788
rect 11032 21732 11036 21788
rect 10972 21728 11036 21732
rect 11052 21788 11116 21792
rect 11052 21732 11056 21788
rect 11056 21732 11112 21788
rect 11112 21732 11116 21788
rect 11052 21728 11116 21732
rect 11132 21788 11196 21792
rect 11132 21732 11136 21788
rect 11136 21732 11192 21788
rect 11192 21732 11196 21788
rect 11132 21728 11196 21732
rect 17079 21788 17143 21792
rect 17079 21732 17083 21788
rect 17083 21732 17139 21788
rect 17139 21732 17143 21788
rect 17079 21728 17143 21732
rect 17159 21788 17223 21792
rect 17159 21732 17163 21788
rect 17163 21732 17219 21788
rect 17219 21732 17223 21788
rect 17159 21728 17223 21732
rect 17239 21788 17303 21792
rect 17239 21732 17243 21788
rect 17243 21732 17299 21788
rect 17299 21732 17303 21788
rect 17239 21728 17303 21732
rect 17319 21788 17383 21792
rect 17319 21732 17323 21788
rect 17323 21732 17379 21788
rect 17379 21732 17383 21788
rect 17319 21728 17383 21732
rect 23266 21788 23330 21792
rect 23266 21732 23270 21788
rect 23270 21732 23326 21788
rect 23326 21732 23330 21788
rect 23266 21728 23330 21732
rect 23346 21788 23410 21792
rect 23346 21732 23350 21788
rect 23350 21732 23406 21788
rect 23406 21732 23410 21788
rect 23346 21728 23410 21732
rect 23426 21788 23490 21792
rect 23426 21732 23430 21788
rect 23430 21732 23486 21788
rect 23486 21732 23490 21788
rect 23426 21728 23490 21732
rect 23506 21788 23570 21792
rect 23506 21732 23510 21788
rect 23510 21732 23566 21788
rect 23566 21732 23570 21788
rect 23506 21728 23570 21732
rect 4045 21244 4109 21248
rect 4045 21188 4049 21244
rect 4049 21188 4105 21244
rect 4105 21188 4109 21244
rect 4045 21184 4109 21188
rect 4125 21244 4189 21248
rect 4125 21188 4129 21244
rect 4129 21188 4185 21244
rect 4185 21188 4189 21244
rect 4125 21184 4189 21188
rect 4205 21244 4269 21248
rect 4205 21188 4209 21244
rect 4209 21188 4265 21244
rect 4265 21188 4269 21244
rect 4205 21184 4269 21188
rect 4285 21244 4349 21248
rect 4285 21188 4289 21244
rect 4289 21188 4345 21244
rect 4345 21188 4349 21244
rect 4285 21184 4349 21188
rect 10232 21244 10296 21248
rect 10232 21188 10236 21244
rect 10236 21188 10292 21244
rect 10292 21188 10296 21244
rect 10232 21184 10296 21188
rect 10312 21244 10376 21248
rect 10312 21188 10316 21244
rect 10316 21188 10372 21244
rect 10372 21188 10376 21244
rect 10312 21184 10376 21188
rect 10392 21244 10456 21248
rect 10392 21188 10396 21244
rect 10396 21188 10452 21244
rect 10452 21188 10456 21244
rect 10392 21184 10456 21188
rect 10472 21244 10536 21248
rect 10472 21188 10476 21244
rect 10476 21188 10532 21244
rect 10532 21188 10536 21244
rect 10472 21184 10536 21188
rect 16419 21244 16483 21248
rect 16419 21188 16423 21244
rect 16423 21188 16479 21244
rect 16479 21188 16483 21244
rect 16419 21184 16483 21188
rect 16499 21244 16563 21248
rect 16499 21188 16503 21244
rect 16503 21188 16559 21244
rect 16559 21188 16563 21244
rect 16499 21184 16563 21188
rect 16579 21244 16643 21248
rect 16579 21188 16583 21244
rect 16583 21188 16639 21244
rect 16639 21188 16643 21244
rect 16579 21184 16643 21188
rect 16659 21244 16723 21248
rect 16659 21188 16663 21244
rect 16663 21188 16719 21244
rect 16719 21188 16723 21244
rect 16659 21184 16723 21188
rect 22606 21244 22670 21248
rect 22606 21188 22610 21244
rect 22610 21188 22666 21244
rect 22666 21188 22670 21244
rect 22606 21184 22670 21188
rect 22686 21244 22750 21248
rect 22686 21188 22690 21244
rect 22690 21188 22746 21244
rect 22746 21188 22750 21244
rect 22686 21184 22750 21188
rect 22766 21244 22830 21248
rect 22766 21188 22770 21244
rect 22770 21188 22826 21244
rect 22826 21188 22830 21244
rect 22766 21184 22830 21188
rect 22846 21244 22910 21248
rect 22846 21188 22850 21244
rect 22850 21188 22906 21244
rect 22906 21188 22910 21244
rect 22846 21184 22910 21188
rect 7788 20768 7852 20772
rect 7788 20712 7838 20768
rect 7838 20712 7852 20768
rect 7788 20708 7852 20712
rect 4705 20700 4769 20704
rect 4705 20644 4709 20700
rect 4709 20644 4765 20700
rect 4765 20644 4769 20700
rect 4705 20640 4769 20644
rect 4785 20700 4849 20704
rect 4785 20644 4789 20700
rect 4789 20644 4845 20700
rect 4845 20644 4849 20700
rect 4785 20640 4849 20644
rect 4865 20700 4929 20704
rect 4865 20644 4869 20700
rect 4869 20644 4925 20700
rect 4925 20644 4929 20700
rect 4865 20640 4929 20644
rect 4945 20700 5009 20704
rect 4945 20644 4949 20700
rect 4949 20644 5005 20700
rect 5005 20644 5009 20700
rect 4945 20640 5009 20644
rect 10892 20700 10956 20704
rect 10892 20644 10896 20700
rect 10896 20644 10952 20700
rect 10952 20644 10956 20700
rect 10892 20640 10956 20644
rect 10972 20700 11036 20704
rect 10972 20644 10976 20700
rect 10976 20644 11032 20700
rect 11032 20644 11036 20700
rect 10972 20640 11036 20644
rect 11052 20700 11116 20704
rect 11052 20644 11056 20700
rect 11056 20644 11112 20700
rect 11112 20644 11116 20700
rect 11052 20640 11116 20644
rect 11132 20700 11196 20704
rect 11132 20644 11136 20700
rect 11136 20644 11192 20700
rect 11192 20644 11196 20700
rect 11132 20640 11196 20644
rect 17079 20700 17143 20704
rect 17079 20644 17083 20700
rect 17083 20644 17139 20700
rect 17139 20644 17143 20700
rect 17079 20640 17143 20644
rect 17159 20700 17223 20704
rect 17159 20644 17163 20700
rect 17163 20644 17219 20700
rect 17219 20644 17223 20700
rect 17159 20640 17223 20644
rect 17239 20700 17303 20704
rect 17239 20644 17243 20700
rect 17243 20644 17299 20700
rect 17299 20644 17303 20700
rect 17239 20640 17303 20644
rect 17319 20700 17383 20704
rect 17319 20644 17323 20700
rect 17323 20644 17379 20700
rect 17379 20644 17383 20700
rect 17319 20640 17383 20644
rect 23266 20700 23330 20704
rect 23266 20644 23270 20700
rect 23270 20644 23326 20700
rect 23326 20644 23330 20700
rect 23266 20640 23330 20644
rect 23346 20700 23410 20704
rect 23346 20644 23350 20700
rect 23350 20644 23406 20700
rect 23406 20644 23410 20700
rect 23346 20640 23410 20644
rect 23426 20700 23490 20704
rect 23426 20644 23430 20700
rect 23430 20644 23486 20700
rect 23486 20644 23490 20700
rect 23426 20640 23490 20644
rect 23506 20700 23570 20704
rect 23506 20644 23510 20700
rect 23510 20644 23566 20700
rect 23566 20644 23570 20700
rect 23506 20640 23570 20644
rect 4045 20156 4109 20160
rect 4045 20100 4049 20156
rect 4049 20100 4105 20156
rect 4105 20100 4109 20156
rect 4045 20096 4109 20100
rect 4125 20156 4189 20160
rect 4125 20100 4129 20156
rect 4129 20100 4185 20156
rect 4185 20100 4189 20156
rect 4125 20096 4189 20100
rect 4205 20156 4269 20160
rect 4205 20100 4209 20156
rect 4209 20100 4265 20156
rect 4265 20100 4269 20156
rect 4205 20096 4269 20100
rect 4285 20156 4349 20160
rect 4285 20100 4289 20156
rect 4289 20100 4345 20156
rect 4345 20100 4349 20156
rect 4285 20096 4349 20100
rect 10232 20156 10296 20160
rect 10232 20100 10236 20156
rect 10236 20100 10292 20156
rect 10292 20100 10296 20156
rect 10232 20096 10296 20100
rect 10312 20156 10376 20160
rect 10312 20100 10316 20156
rect 10316 20100 10372 20156
rect 10372 20100 10376 20156
rect 10312 20096 10376 20100
rect 10392 20156 10456 20160
rect 10392 20100 10396 20156
rect 10396 20100 10452 20156
rect 10452 20100 10456 20156
rect 10392 20096 10456 20100
rect 10472 20156 10536 20160
rect 10472 20100 10476 20156
rect 10476 20100 10532 20156
rect 10532 20100 10536 20156
rect 10472 20096 10536 20100
rect 16419 20156 16483 20160
rect 16419 20100 16423 20156
rect 16423 20100 16479 20156
rect 16479 20100 16483 20156
rect 16419 20096 16483 20100
rect 16499 20156 16563 20160
rect 16499 20100 16503 20156
rect 16503 20100 16559 20156
rect 16559 20100 16563 20156
rect 16499 20096 16563 20100
rect 16579 20156 16643 20160
rect 16579 20100 16583 20156
rect 16583 20100 16639 20156
rect 16639 20100 16643 20156
rect 16579 20096 16643 20100
rect 16659 20156 16723 20160
rect 16659 20100 16663 20156
rect 16663 20100 16719 20156
rect 16719 20100 16723 20156
rect 16659 20096 16723 20100
rect 22606 20156 22670 20160
rect 22606 20100 22610 20156
rect 22610 20100 22666 20156
rect 22666 20100 22670 20156
rect 22606 20096 22670 20100
rect 22686 20156 22750 20160
rect 22686 20100 22690 20156
rect 22690 20100 22746 20156
rect 22746 20100 22750 20156
rect 22686 20096 22750 20100
rect 22766 20156 22830 20160
rect 22766 20100 22770 20156
rect 22770 20100 22826 20156
rect 22826 20100 22830 20156
rect 22766 20096 22830 20100
rect 22846 20156 22910 20160
rect 22846 20100 22850 20156
rect 22850 20100 22906 20156
rect 22906 20100 22910 20156
rect 22846 20096 22910 20100
rect 4705 19612 4769 19616
rect 4705 19556 4709 19612
rect 4709 19556 4765 19612
rect 4765 19556 4769 19612
rect 4705 19552 4769 19556
rect 4785 19612 4849 19616
rect 4785 19556 4789 19612
rect 4789 19556 4845 19612
rect 4845 19556 4849 19612
rect 4785 19552 4849 19556
rect 4865 19612 4929 19616
rect 4865 19556 4869 19612
rect 4869 19556 4925 19612
rect 4925 19556 4929 19612
rect 4865 19552 4929 19556
rect 4945 19612 5009 19616
rect 4945 19556 4949 19612
rect 4949 19556 5005 19612
rect 5005 19556 5009 19612
rect 4945 19552 5009 19556
rect 10892 19612 10956 19616
rect 10892 19556 10896 19612
rect 10896 19556 10952 19612
rect 10952 19556 10956 19612
rect 10892 19552 10956 19556
rect 10972 19612 11036 19616
rect 10972 19556 10976 19612
rect 10976 19556 11032 19612
rect 11032 19556 11036 19612
rect 10972 19552 11036 19556
rect 11052 19612 11116 19616
rect 11052 19556 11056 19612
rect 11056 19556 11112 19612
rect 11112 19556 11116 19612
rect 11052 19552 11116 19556
rect 11132 19612 11196 19616
rect 11132 19556 11136 19612
rect 11136 19556 11192 19612
rect 11192 19556 11196 19612
rect 11132 19552 11196 19556
rect 17079 19612 17143 19616
rect 17079 19556 17083 19612
rect 17083 19556 17139 19612
rect 17139 19556 17143 19612
rect 17079 19552 17143 19556
rect 17159 19612 17223 19616
rect 17159 19556 17163 19612
rect 17163 19556 17219 19612
rect 17219 19556 17223 19612
rect 17159 19552 17223 19556
rect 17239 19612 17303 19616
rect 17239 19556 17243 19612
rect 17243 19556 17299 19612
rect 17299 19556 17303 19612
rect 17239 19552 17303 19556
rect 17319 19612 17383 19616
rect 17319 19556 17323 19612
rect 17323 19556 17379 19612
rect 17379 19556 17383 19612
rect 17319 19552 17383 19556
rect 23266 19612 23330 19616
rect 23266 19556 23270 19612
rect 23270 19556 23326 19612
rect 23326 19556 23330 19612
rect 23266 19552 23330 19556
rect 23346 19612 23410 19616
rect 23346 19556 23350 19612
rect 23350 19556 23406 19612
rect 23406 19556 23410 19612
rect 23346 19552 23410 19556
rect 23426 19612 23490 19616
rect 23426 19556 23430 19612
rect 23430 19556 23486 19612
rect 23486 19556 23490 19612
rect 23426 19552 23490 19556
rect 23506 19612 23570 19616
rect 23506 19556 23510 19612
rect 23510 19556 23566 19612
rect 23566 19556 23570 19612
rect 23506 19552 23570 19556
rect 4045 19068 4109 19072
rect 4045 19012 4049 19068
rect 4049 19012 4105 19068
rect 4105 19012 4109 19068
rect 4045 19008 4109 19012
rect 4125 19068 4189 19072
rect 4125 19012 4129 19068
rect 4129 19012 4185 19068
rect 4185 19012 4189 19068
rect 4125 19008 4189 19012
rect 4205 19068 4269 19072
rect 4205 19012 4209 19068
rect 4209 19012 4265 19068
rect 4265 19012 4269 19068
rect 4205 19008 4269 19012
rect 4285 19068 4349 19072
rect 4285 19012 4289 19068
rect 4289 19012 4345 19068
rect 4345 19012 4349 19068
rect 4285 19008 4349 19012
rect 10232 19068 10296 19072
rect 10232 19012 10236 19068
rect 10236 19012 10292 19068
rect 10292 19012 10296 19068
rect 10232 19008 10296 19012
rect 10312 19068 10376 19072
rect 10312 19012 10316 19068
rect 10316 19012 10372 19068
rect 10372 19012 10376 19068
rect 10312 19008 10376 19012
rect 10392 19068 10456 19072
rect 10392 19012 10396 19068
rect 10396 19012 10452 19068
rect 10452 19012 10456 19068
rect 10392 19008 10456 19012
rect 10472 19068 10536 19072
rect 10472 19012 10476 19068
rect 10476 19012 10532 19068
rect 10532 19012 10536 19068
rect 10472 19008 10536 19012
rect 16419 19068 16483 19072
rect 16419 19012 16423 19068
rect 16423 19012 16479 19068
rect 16479 19012 16483 19068
rect 16419 19008 16483 19012
rect 16499 19068 16563 19072
rect 16499 19012 16503 19068
rect 16503 19012 16559 19068
rect 16559 19012 16563 19068
rect 16499 19008 16563 19012
rect 16579 19068 16643 19072
rect 16579 19012 16583 19068
rect 16583 19012 16639 19068
rect 16639 19012 16643 19068
rect 16579 19008 16643 19012
rect 16659 19068 16723 19072
rect 16659 19012 16663 19068
rect 16663 19012 16719 19068
rect 16719 19012 16723 19068
rect 16659 19008 16723 19012
rect 22606 19068 22670 19072
rect 22606 19012 22610 19068
rect 22610 19012 22666 19068
rect 22666 19012 22670 19068
rect 22606 19008 22670 19012
rect 22686 19068 22750 19072
rect 22686 19012 22690 19068
rect 22690 19012 22746 19068
rect 22746 19012 22750 19068
rect 22686 19008 22750 19012
rect 22766 19068 22830 19072
rect 22766 19012 22770 19068
rect 22770 19012 22826 19068
rect 22826 19012 22830 19068
rect 22766 19008 22830 19012
rect 22846 19068 22910 19072
rect 22846 19012 22850 19068
rect 22850 19012 22906 19068
rect 22906 19012 22910 19068
rect 22846 19008 22910 19012
rect 4705 18524 4769 18528
rect 4705 18468 4709 18524
rect 4709 18468 4765 18524
rect 4765 18468 4769 18524
rect 4705 18464 4769 18468
rect 4785 18524 4849 18528
rect 4785 18468 4789 18524
rect 4789 18468 4845 18524
rect 4845 18468 4849 18524
rect 4785 18464 4849 18468
rect 4865 18524 4929 18528
rect 4865 18468 4869 18524
rect 4869 18468 4925 18524
rect 4925 18468 4929 18524
rect 4865 18464 4929 18468
rect 4945 18524 5009 18528
rect 4945 18468 4949 18524
rect 4949 18468 5005 18524
rect 5005 18468 5009 18524
rect 4945 18464 5009 18468
rect 10892 18524 10956 18528
rect 10892 18468 10896 18524
rect 10896 18468 10952 18524
rect 10952 18468 10956 18524
rect 10892 18464 10956 18468
rect 10972 18524 11036 18528
rect 10972 18468 10976 18524
rect 10976 18468 11032 18524
rect 11032 18468 11036 18524
rect 10972 18464 11036 18468
rect 11052 18524 11116 18528
rect 11052 18468 11056 18524
rect 11056 18468 11112 18524
rect 11112 18468 11116 18524
rect 11052 18464 11116 18468
rect 11132 18524 11196 18528
rect 11132 18468 11136 18524
rect 11136 18468 11192 18524
rect 11192 18468 11196 18524
rect 11132 18464 11196 18468
rect 17079 18524 17143 18528
rect 17079 18468 17083 18524
rect 17083 18468 17139 18524
rect 17139 18468 17143 18524
rect 17079 18464 17143 18468
rect 17159 18524 17223 18528
rect 17159 18468 17163 18524
rect 17163 18468 17219 18524
rect 17219 18468 17223 18524
rect 17159 18464 17223 18468
rect 17239 18524 17303 18528
rect 17239 18468 17243 18524
rect 17243 18468 17299 18524
rect 17299 18468 17303 18524
rect 17239 18464 17303 18468
rect 17319 18524 17383 18528
rect 17319 18468 17323 18524
rect 17323 18468 17379 18524
rect 17379 18468 17383 18524
rect 17319 18464 17383 18468
rect 23266 18524 23330 18528
rect 23266 18468 23270 18524
rect 23270 18468 23326 18524
rect 23326 18468 23330 18524
rect 23266 18464 23330 18468
rect 23346 18524 23410 18528
rect 23346 18468 23350 18524
rect 23350 18468 23406 18524
rect 23406 18468 23410 18524
rect 23346 18464 23410 18468
rect 23426 18524 23490 18528
rect 23426 18468 23430 18524
rect 23430 18468 23486 18524
rect 23486 18468 23490 18524
rect 23426 18464 23490 18468
rect 23506 18524 23570 18528
rect 23506 18468 23510 18524
rect 23510 18468 23566 18524
rect 23566 18468 23570 18524
rect 23506 18464 23570 18468
rect 4045 17980 4109 17984
rect 4045 17924 4049 17980
rect 4049 17924 4105 17980
rect 4105 17924 4109 17980
rect 4045 17920 4109 17924
rect 4125 17980 4189 17984
rect 4125 17924 4129 17980
rect 4129 17924 4185 17980
rect 4185 17924 4189 17980
rect 4125 17920 4189 17924
rect 4205 17980 4269 17984
rect 4205 17924 4209 17980
rect 4209 17924 4265 17980
rect 4265 17924 4269 17980
rect 4205 17920 4269 17924
rect 4285 17980 4349 17984
rect 4285 17924 4289 17980
rect 4289 17924 4345 17980
rect 4345 17924 4349 17980
rect 4285 17920 4349 17924
rect 10232 17980 10296 17984
rect 10232 17924 10236 17980
rect 10236 17924 10292 17980
rect 10292 17924 10296 17980
rect 10232 17920 10296 17924
rect 10312 17980 10376 17984
rect 10312 17924 10316 17980
rect 10316 17924 10372 17980
rect 10372 17924 10376 17980
rect 10312 17920 10376 17924
rect 10392 17980 10456 17984
rect 10392 17924 10396 17980
rect 10396 17924 10452 17980
rect 10452 17924 10456 17980
rect 10392 17920 10456 17924
rect 10472 17980 10536 17984
rect 10472 17924 10476 17980
rect 10476 17924 10532 17980
rect 10532 17924 10536 17980
rect 10472 17920 10536 17924
rect 16419 17980 16483 17984
rect 16419 17924 16423 17980
rect 16423 17924 16479 17980
rect 16479 17924 16483 17980
rect 16419 17920 16483 17924
rect 16499 17980 16563 17984
rect 16499 17924 16503 17980
rect 16503 17924 16559 17980
rect 16559 17924 16563 17980
rect 16499 17920 16563 17924
rect 16579 17980 16643 17984
rect 16579 17924 16583 17980
rect 16583 17924 16639 17980
rect 16639 17924 16643 17980
rect 16579 17920 16643 17924
rect 16659 17980 16723 17984
rect 16659 17924 16663 17980
rect 16663 17924 16719 17980
rect 16719 17924 16723 17980
rect 16659 17920 16723 17924
rect 22606 17980 22670 17984
rect 22606 17924 22610 17980
rect 22610 17924 22666 17980
rect 22666 17924 22670 17980
rect 22606 17920 22670 17924
rect 22686 17980 22750 17984
rect 22686 17924 22690 17980
rect 22690 17924 22746 17980
rect 22746 17924 22750 17980
rect 22686 17920 22750 17924
rect 22766 17980 22830 17984
rect 22766 17924 22770 17980
rect 22770 17924 22826 17980
rect 22826 17924 22830 17980
rect 22766 17920 22830 17924
rect 22846 17980 22910 17984
rect 22846 17924 22850 17980
rect 22850 17924 22906 17980
rect 22906 17924 22910 17980
rect 22846 17920 22910 17924
rect 7788 17852 7852 17916
rect 4705 17436 4769 17440
rect 4705 17380 4709 17436
rect 4709 17380 4765 17436
rect 4765 17380 4769 17436
rect 4705 17376 4769 17380
rect 4785 17436 4849 17440
rect 4785 17380 4789 17436
rect 4789 17380 4845 17436
rect 4845 17380 4849 17436
rect 4785 17376 4849 17380
rect 4865 17436 4929 17440
rect 4865 17380 4869 17436
rect 4869 17380 4925 17436
rect 4925 17380 4929 17436
rect 4865 17376 4929 17380
rect 4945 17436 5009 17440
rect 4945 17380 4949 17436
rect 4949 17380 5005 17436
rect 5005 17380 5009 17436
rect 4945 17376 5009 17380
rect 10892 17436 10956 17440
rect 10892 17380 10896 17436
rect 10896 17380 10952 17436
rect 10952 17380 10956 17436
rect 10892 17376 10956 17380
rect 10972 17436 11036 17440
rect 10972 17380 10976 17436
rect 10976 17380 11032 17436
rect 11032 17380 11036 17436
rect 10972 17376 11036 17380
rect 11052 17436 11116 17440
rect 11052 17380 11056 17436
rect 11056 17380 11112 17436
rect 11112 17380 11116 17436
rect 11052 17376 11116 17380
rect 11132 17436 11196 17440
rect 11132 17380 11136 17436
rect 11136 17380 11192 17436
rect 11192 17380 11196 17436
rect 11132 17376 11196 17380
rect 17079 17436 17143 17440
rect 17079 17380 17083 17436
rect 17083 17380 17139 17436
rect 17139 17380 17143 17436
rect 17079 17376 17143 17380
rect 17159 17436 17223 17440
rect 17159 17380 17163 17436
rect 17163 17380 17219 17436
rect 17219 17380 17223 17436
rect 17159 17376 17223 17380
rect 17239 17436 17303 17440
rect 17239 17380 17243 17436
rect 17243 17380 17299 17436
rect 17299 17380 17303 17436
rect 17239 17376 17303 17380
rect 17319 17436 17383 17440
rect 17319 17380 17323 17436
rect 17323 17380 17379 17436
rect 17379 17380 17383 17436
rect 17319 17376 17383 17380
rect 23266 17436 23330 17440
rect 23266 17380 23270 17436
rect 23270 17380 23326 17436
rect 23326 17380 23330 17436
rect 23266 17376 23330 17380
rect 23346 17436 23410 17440
rect 23346 17380 23350 17436
rect 23350 17380 23406 17436
rect 23406 17380 23410 17436
rect 23346 17376 23410 17380
rect 23426 17436 23490 17440
rect 23426 17380 23430 17436
rect 23430 17380 23486 17436
rect 23486 17380 23490 17436
rect 23426 17376 23490 17380
rect 23506 17436 23570 17440
rect 23506 17380 23510 17436
rect 23510 17380 23566 17436
rect 23566 17380 23570 17436
rect 23506 17376 23570 17380
rect 4045 16892 4109 16896
rect 4045 16836 4049 16892
rect 4049 16836 4105 16892
rect 4105 16836 4109 16892
rect 4045 16832 4109 16836
rect 4125 16892 4189 16896
rect 4125 16836 4129 16892
rect 4129 16836 4185 16892
rect 4185 16836 4189 16892
rect 4125 16832 4189 16836
rect 4205 16892 4269 16896
rect 4205 16836 4209 16892
rect 4209 16836 4265 16892
rect 4265 16836 4269 16892
rect 4205 16832 4269 16836
rect 4285 16892 4349 16896
rect 4285 16836 4289 16892
rect 4289 16836 4345 16892
rect 4345 16836 4349 16892
rect 4285 16832 4349 16836
rect 10232 16892 10296 16896
rect 10232 16836 10236 16892
rect 10236 16836 10292 16892
rect 10292 16836 10296 16892
rect 10232 16832 10296 16836
rect 10312 16892 10376 16896
rect 10312 16836 10316 16892
rect 10316 16836 10372 16892
rect 10372 16836 10376 16892
rect 10312 16832 10376 16836
rect 10392 16892 10456 16896
rect 10392 16836 10396 16892
rect 10396 16836 10452 16892
rect 10452 16836 10456 16892
rect 10392 16832 10456 16836
rect 10472 16892 10536 16896
rect 10472 16836 10476 16892
rect 10476 16836 10532 16892
rect 10532 16836 10536 16892
rect 10472 16832 10536 16836
rect 16419 16892 16483 16896
rect 16419 16836 16423 16892
rect 16423 16836 16479 16892
rect 16479 16836 16483 16892
rect 16419 16832 16483 16836
rect 16499 16892 16563 16896
rect 16499 16836 16503 16892
rect 16503 16836 16559 16892
rect 16559 16836 16563 16892
rect 16499 16832 16563 16836
rect 16579 16892 16643 16896
rect 16579 16836 16583 16892
rect 16583 16836 16639 16892
rect 16639 16836 16643 16892
rect 16579 16832 16643 16836
rect 16659 16892 16723 16896
rect 16659 16836 16663 16892
rect 16663 16836 16719 16892
rect 16719 16836 16723 16892
rect 16659 16832 16723 16836
rect 22606 16892 22670 16896
rect 22606 16836 22610 16892
rect 22610 16836 22666 16892
rect 22666 16836 22670 16892
rect 22606 16832 22670 16836
rect 22686 16892 22750 16896
rect 22686 16836 22690 16892
rect 22690 16836 22746 16892
rect 22746 16836 22750 16892
rect 22686 16832 22750 16836
rect 22766 16892 22830 16896
rect 22766 16836 22770 16892
rect 22770 16836 22826 16892
rect 22826 16836 22830 16892
rect 22766 16832 22830 16836
rect 22846 16892 22910 16896
rect 22846 16836 22850 16892
rect 22850 16836 22906 16892
rect 22906 16836 22910 16892
rect 22846 16832 22910 16836
rect 4705 16348 4769 16352
rect 4705 16292 4709 16348
rect 4709 16292 4765 16348
rect 4765 16292 4769 16348
rect 4705 16288 4769 16292
rect 4785 16348 4849 16352
rect 4785 16292 4789 16348
rect 4789 16292 4845 16348
rect 4845 16292 4849 16348
rect 4785 16288 4849 16292
rect 4865 16348 4929 16352
rect 4865 16292 4869 16348
rect 4869 16292 4925 16348
rect 4925 16292 4929 16348
rect 4865 16288 4929 16292
rect 4945 16348 5009 16352
rect 4945 16292 4949 16348
rect 4949 16292 5005 16348
rect 5005 16292 5009 16348
rect 4945 16288 5009 16292
rect 10892 16348 10956 16352
rect 10892 16292 10896 16348
rect 10896 16292 10952 16348
rect 10952 16292 10956 16348
rect 10892 16288 10956 16292
rect 10972 16348 11036 16352
rect 10972 16292 10976 16348
rect 10976 16292 11032 16348
rect 11032 16292 11036 16348
rect 10972 16288 11036 16292
rect 11052 16348 11116 16352
rect 11052 16292 11056 16348
rect 11056 16292 11112 16348
rect 11112 16292 11116 16348
rect 11052 16288 11116 16292
rect 11132 16348 11196 16352
rect 11132 16292 11136 16348
rect 11136 16292 11192 16348
rect 11192 16292 11196 16348
rect 11132 16288 11196 16292
rect 17079 16348 17143 16352
rect 17079 16292 17083 16348
rect 17083 16292 17139 16348
rect 17139 16292 17143 16348
rect 17079 16288 17143 16292
rect 17159 16348 17223 16352
rect 17159 16292 17163 16348
rect 17163 16292 17219 16348
rect 17219 16292 17223 16348
rect 17159 16288 17223 16292
rect 17239 16348 17303 16352
rect 17239 16292 17243 16348
rect 17243 16292 17299 16348
rect 17299 16292 17303 16348
rect 17239 16288 17303 16292
rect 17319 16348 17383 16352
rect 17319 16292 17323 16348
rect 17323 16292 17379 16348
rect 17379 16292 17383 16348
rect 17319 16288 17383 16292
rect 23266 16348 23330 16352
rect 23266 16292 23270 16348
rect 23270 16292 23326 16348
rect 23326 16292 23330 16348
rect 23266 16288 23330 16292
rect 23346 16348 23410 16352
rect 23346 16292 23350 16348
rect 23350 16292 23406 16348
rect 23406 16292 23410 16348
rect 23346 16288 23410 16292
rect 23426 16348 23490 16352
rect 23426 16292 23430 16348
rect 23430 16292 23486 16348
rect 23486 16292 23490 16348
rect 23426 16288 23490 16292
rect 23506 16348 23570 16352
rect 23506 16292 23510 16348
rect 23510 16292 23566 16348
rect 23566 16292 23570 16348
rect 23506 16288 23570 16292
rect 4045 15804 4109 15808
rect 4045 15748 4049 15804
rect 4049 15748 4105 15804
rect 4105 15748 4109 15804
rect 4045 15744 4109 15748
rect 4125 15804 4189 15808
rect 4125 15748 4129 15804
rect 4129 15748 4185 15804
rect 4185 15748 4189 15804
rect 4125 15744 4189 15748
rect 4205 15804 4269 15808
rect 4205 15748 4209 15804
rect 4209 15748 4265 15804
rect 4265 15748 4269 15804
rect 4205 15744 4269 15748
rect 4285 15804 4349 15808
rect 4285 15748 4289 15804
rect 4289 15748 4345 15804
rect 4345 15748 4349 15804
rect 4285 15744 4349 15748
rect 10232 15804 10296 15808
rect 10232 15748 10236 15804
rect 10236 15748 10292 15804
rect 10292 15748 10296 15804
rect 10232 15744 10296 15748
rect 10312 15804 10376 15808
rect 10312 15748 10316 15804
rect 10316 15748 10372 15804
rect 10372 15748 10376 15804
rect 10312 15744 10376 15748
rect 10392 15804 10456 15808
rect 10392 15748 10396 15804
rect 10396 15748 10452 15804
rect 10452 15748 10456 15804
rect 10392 15744 10456 15748
rect 10472 15804 10536 15808
rect 10472 15748 10476 15804
rect 10476 15748 10532 15804
rect 10532 15748 10536 15804
rect 10472 15744 10536 15748
rect 16419 15804 16483 15808
rect 16419 15748 16423 15804
rect 16423 15748 16479 15804
rect 16479 15748 16483 15804
rect 16419 15744 16483 15748
rect 16499 15804 16563 15808
rect 16499 15748 16503 15804
rect 16503 15748 16559 15804
rect 16559 15748 16563 15804
rect 16499 15744 16563 15748
rect 16579 15804 16643 15808
rect 16579 15748 16583 15804
rect 16583 15748 16639 15804
rect 16639 15748 16643 15804
rect 16579 15744 16643 15748
rect 16659 15804 16723 15808
rect 16659 15748 16663 15804
rect 16663 15748 16719 15804
rect 16719 15748 16723 15804
rect 16659 15744 16723 15748
rect 22606 15804 22670 15808
rect 22606 15748 22610 15804
rect 22610 15748 22666 15804
rect 22666 15748 22670 15804
rect 22606 15744 22670 15748
rect 22686 15804 22750 15808
rect 22686 15748 22690 15804
rect 22690 15748 22746 15804
rect 22746 15748 22750 15804
rect 22686 15744 22750 15748
rect 22766 15804 22830 15808
rect 22766 15748 22770 15804
rect 22770 15748 22826 15804
rect 22826 15748 22830 15804
rect 22766 15744 22830 15748
rect 22846 15804 22910 15808
rect 22846 15748 22850 15804
rect 22850 15748 22906 15804
rect 22906 15748 22910 15804
rect 22846 15744 22910 15748
rect 4705 15260 4769 15264
rect 4705 15204 4709 15260
rect 4709 15204 4765 15260
rect 4765 15204 4769 15260
rect 4705 15200 4769 15204
rect 4785 15260 4849 15264
rect 4785 15204 4789 15260
rect 4789 15204 4845 15260
rect 4845 15204 4849 15260
rect 4785 15200 4849 15204
rect 4865 15260 4929 15264
rect 4865 15204 4869 15260
rect 4869 15204 4925 15260
rect 4925 15204 4929 15260
rect 4865 15200 4929 15204
rect 4945 15260 5009 15264
rect 4945 15204 4949 15260
rect 4949 15204 5005 15260
rect 5005 15204 5009 15260
rect 4945 15200 5009 15204
rect 10892 15260 10956 15264
rect 10892 15204 10896 15260
rect 10896 15204 10952 15260
rect 10952 15204 10956 15260
rect 10892 15200 10956 15204
rect 10972 15260 11036 15264
rect 10972 15204 10976 15260
rect 10976 15204 11032 15260
rect 11032 15204 11036 15260
rect 10972 15200 11036 15204
rect 11052 15260 11116 15264
rect 11052 15204 11056 15260
rect 11056 15204 11112 15260
rect 11112 15204 11116 15260
rect 11052 15200 11116 15204
rect 11132 15260 11196 15264
rect 11132 15204 11136 15260
rect 11136 15204 11192 15260
rect 11192 15204 11196 15260
rect 11132 15200 11196 15204
rect 17079 15260 17143 15264
rect 17079 15204 17083 15260
rect 17083 15204 17139 15260
rect 17139 15204 17143 15260
rect 17079 15200 17143 15204
rect 17159 15260 17223 15264
rect 17159 15204 17163 15260
rect 17163 15204 17219 15260
rect 17219 15204 17223 15260
rect 17159 15200 17223 15204
rect 17239 15260 17303 15264
rect 17239 15204 17243 15260
rect 17243 15204 17299 15260
rect 17299 15204 17303 15260
rect 17239 15200 17303 15204
rect 17319 15260 17383 15264
rect 17319 15204 17323 15260
rect 17323 15204 17379 15260
rect 17379 15204 17383 15260
rect 17319 15200 17383 15204
rect 23266 15260 23330 15264
rect 23266 15204 23270 15260
rect 23270 15204 23326 15260
rect 23326 15204 23330 15260
rect 23266 15200 23330 15204
rect 23346 15260 23410 15264
rect 23346 15204 23350 15260
rect 23350 15204 23406 15260
rect 23406 15204 23410 15260
rect 23346 15200 23410 15204
rect 23426 15260 23490 15264
rect 23426 15204 23430 15260
rect 23430 15204 23486 15260
rect 23486 15204 23490 15260
rect 23426 15200 23490 15204
rect 23506 15260 23570 15264
rect 23506 15204 23510 15260
rect 23510 15204 23566 15260
rect 23566 15204 23570 15260
rect 23506 15200 23570 15204
rect 4045 14716 4109 14720
rect 4045 14660 4049 14716
rect 4049 14660 4105 14716
rect 4105 14660 4109 14716
rect 4045 14656 4109 14660
rect 4125 14716 4189 14720
rect 4125 14660 4129 14716
rect 4129 14660 4185 14716
rect 4185 14660 4189 14716
rect 4125 14656 4189 14660
rect 4205 14716 4269 14720
rect 4205 14660 4209 14716
rect 4209 14660 4265 14716
rect 4265 14660 4269 14716
rect 4205 14656 4269 14660
rect 4285 14716 4349 14720
rect 4285 14660 4289 14716
rect 4289 14660 4345 14716
rect 4345 14660 4349 14716
rect 4285 14656 4349 14660
rect 10232 14716 10296 14720
rect 10232 14660 10236 14716
rect 10236 14660 10292 14716
rect 10292 14660 10296 14716
rect 10232 14656 10296 14660
rect 10312 14716 10376 14720
rect 10312 14660 10316 14716
rect 10316 14660 10372 14716
rect 10372 14660 10376 14716
rect 10312 14656 10376 14660
rect 10392 14716 10456 14720
rect 10392 14660 10396 14716
rect 10396 14660 10452 14716
rect 10452 14660 10456 14716
rect 10392 14656 10456 14660
rect 10472 14716 10536 14720
rect 10472 14660 10476 14716
rect 10476 14660 10532 14716
rect 10532 14660 10536 14716
rect 10472 14656 10536 14660
rect 16419 14716 16483 14720
rect 16419 14660 16423 14716
rect 16423 14660 16479 14716
rect 16479 14660 16483 14716
rect 16419 14656 16483 14660
rect 16499 14716 16563 14720
rect 16499 14660 16503 14716
rect 16503 14660 16559 14716
rect 16559 14660 16563 14716
rect 16499 14656 16563 14660
rect 16579 14716 16643 14720
rect 16579 14660 16583 14716
rect 16583 14660 16639 14716
rect 16639 14660 16643 14716
rect 16579 14656 16643 14660
rect 16659 14716 16723 14720
rect 16659 14660 16663 14716
rect 16663 14660 16719 14716
rect 16719 14660 16723 14716
rect 16659 14656 16723 14660
rect 22606 14716 22670 14720
rect 22606 14660 22610 14716
rect 22610 14660 22666 14716
rect 22666 14660 22670 14716
rect 22606 14656 22670 14660
rect 22686 14716 22750 14720
rect 22686 14660 22690 14716
rect 22690 14660 22746 14716
rect 22746 14660 22750 14716
rect 22686 14656 22750 14660
rect 22766 14716 22830 14720
rect 22766 14660 22770 14716
rect 22770 14660 22826 14716
rect 22826 14660 22830 14716
rect 22766 14656 22830 14660
rect 22846 14716 22910 14720
rect 22846 14660 22850 14716
rect 22850 14660 22906 14716
rect 22906 14660 22910 14716
rect 22846 14656 22910 14660
rect 4705 14172 4769 14176
rect 4705 14116 4709 14172
rect 4709 14116 4765 14172
rect 4765 14116 4769 14172
rect 4705 14112 4769 14116
rect 4785 14172 4849 14176
rect 4785 14116 4789 14172
rect 4789 14116 4845 14172
rect 4845 14116 4849 14172
rect 4785 14112 4849 14116
rect 4865 14172 4929 14176
rect 4865 14116 4869 14172
rect 4869 14116 4925 14172
rect 4925 14116 4929 14172
rect 4865 14112 4929 14116
rect 4945 14172 5009 14176
rect 4945 14116 4949 14172
rect 4949 14116 5005 14172
rect 5005 14116 5009 14172
rect 4945 14112 5009 14116
rect 10892 14172 10956 14176
rect 10892 14116 10896 14172
rect 10896 14116 10952 14172
rect 10952 14116 10956 14172
rect 10892 14112 10956 14116
rect 10972 14172 11036 14176
rect 10972 14116 10976 14172
rect 10976 14116 11032 14172
rect 11032 14116 11036 14172
rect 10972 14112 11036 14116
rect 11052 14172 11116 14176
rect 11052 14116 11056 14172
rect 11056 14116 11112 14172
rect 11112 14116 11116 14172
rect 11052 14112 11116 14116
rect 11132 14172 11196 14176
rect 11132 14116 11136 14172
rect 11136 14116 11192 14172
rect 11192 14116 11196 14172
rect 11132 14112 11196 14116
rect 17079 14172 17143 14176
rect 17079 14116 17083 14172
rect 17083 14116 17139 14172
rect 17139 14116 17143 14172
rect 17079 14112 17143 14116
rect 17159 14172 17223 14176
rect 17159 14116 17163 14172
rect 17163 14116 17219 14172
rect 17219 14116 17223 14172
rect 17159 14112 17223 14116
rect 17239 14172 17303 14176
rect 17239 14116 17243 14172
rect 17243 14116 17299 14172
rect 17299 14116 17303 14172
rect 17239 14112 17303 14116
rect 17319 14172 17383 14176
rect 17319 14116 17323 14172
rect 17323 14116 17379 14172
rect 17379 14116 17383 14172
rect 17319 14112 17383 14116
rect 23266 14172 23330 14176
rect 23266 14116 23270 14172
rect 23270 14116 23326 14172
rect 23326 14116 23330 14172
rect 23266 14112 23330 14116
rect 23346 14172 23410 14176
rect 23346 14116 23350 14172
rect 23350 14116 23406 14172
rect 23406 14116 23410 14172
rect 23346 14112 23410 14116
rect 23426 14172 23490 14176
rect 23426 14116 23430 14172
rect 23430 14116 23486 14172
rect 23486 14116 23490 14172
rect 23426 14112 23490 14116
rect 23506 14172 23570 14176
rect 23506 14116 23510 14172
rect 23510 14116 23566 14172
rect 23566 14116 23570 14172
rect 23506 14112 23570 14116
rect 4045 13628 4109 13632
rect 4045 13572 4049 13628
rect 4049 13572 4105 13628
rect 4105 13572 4109 13628
rect 4045 13568 4109 13572
rect 4125 13628 4189 13632
rect 4125 13572 4129 13628
rect 4129 13572 4185 13628
rect 4185 13572 4189 13628
rect 4125 13568 4189 13572
rect 4205 13628 4269 13632
rect 4205 13572 4209 13628
rect 4209 13572 4265 13628
rect 4265 13572 4269 13628
rect 4205 13568 4269 13572
rect 4285 13628 4349 13632
rect 4285 13572 4289 13628
rect 4289 13572 4345 13628
rect 4345 13572 4349 13628
rect 4285 13568 4349 13572
rect 10232 13628 10296 13632
rect 10232 13572 10236 13628
rect 10236 13572 10292 13628
rect 10292 13572 10296 13628
rect 10232 13568 10296 13572
rect 10312 13628 10376 13632
rect 10312 13572 10316 13628
rect 10316 13572 10372 13628
rect 10372 13572 10376 13628
rect 10312 13568 10376 13572
rect 10392 13628 10456 13632
rect 10392 13572 10396 13628
rect 10396 13572 10452 13628
rect 10452 13572 10456 13628
rect 10392 13568 10456 13572
rect 10472 13628 10536 13632
rect 10472 13572 10476 13628
rect 10476 13572 10532 13628
rect 10532 13572 10536 13628
rect 10472 13568 10536 13572
rect 16419 13628 16483 13632
rect 16419 13572 16423 13628
rect 16423 13572 16479 13628
rect 16479 13572 16483 13628
rect 16419 13568 16483 13572
rect 16499 13628 16563 13632
rect 16499 13572 16503 13628
rect 16503 13572 16559 13628
rect 16559 13572 16563 13628
rect 16499 13568 16563 13572
rect 16579 13628 16643 13632
rect 16579 13572 16583 13628
rect 16583 13572 16639 13628
rect 16639 13572 16643 13628
rect 16579 13568 16643 13572
rect 16659 13628 16723 13632
rect 16659 13572 16663 13628
rect 16663 13572 16719 13628
rect 16719 13572 16723 13628
rect 16659 13568 16723 13572
rect 22606 13628 22670 13632
rect 22606 13572 22610 13628
rect 22610 13572 22666 13628
rect 22666 13572 22670 13628
rect 22606 13568 22670 13572
rect 22686 13628 22750 13632
rect 22686 13572 22690 13628
rect 22690 13572 22746 13628
rect 22746 13572 22750 13628
rect 22686 13568 22750 13572
rect 22766 13628 22830 13632
rect 22766 13572 22770 13628
rect 22770 13572 22826 13628
rect 22826 13572 22830 13628
rect 22766 13568 22830 13572
rect 22846 13628 22910 13632
rect 22846 13572 22850 13628
rect 22850 13572 22906 13628
rect 22906 13572 22910 13628
rect 22846 13568 22910 13572
rect 4705 13084 4769 13088
rect 4705 13028 4709 13084
rect 4709 13028 4765 13084
rect 4765 13028 4769 13084
rect 4705 13024 4769 13028
rect 4785 13084 4849 13088
rect 4785 13028 4789 13084
rect 4789 13028 4845 13084
rect 4845 13028 4849 13084
rect 4785 13024 4849 13028
rect 4865 13084 4929 13088
rect 4865 13028 4869 13084
rect 4869 13028 4925 13084
rect 4925 13028 4929 13084
rect 4865 13024 4929 13028
rect 4945 13084 5009 13088
rect 4945 13028 4949 13084
rect 4949 13028 5005 13084
rect 5005 13028 5009 13084
rect 4945 13024 5009 13028
rect 10892 13084 10956 13088
rect 10892 13028 10896 13084
rect 10896 13028 10952 13084
rect 10952 13028 10956 13084
rect 10892 13024 10956 13028
rect 10972 13084 11036 13088
rect 10972 13028 10976 13084
rect 10976 13028 11032 13084
rect 11032 13028 11036 13084
rect 10972 13024 11036 13028
rect 11052 13084 11116 13088
rect 11052 13028 11056 13084
rect 11056 13028 11112 13084
rect 11112 13028 11116 13084
rect 11052 13024 11116 13028
rect 11132 13084 11196 13088
rect 11132 13028 11136 13084
rect 11136 13028 11192 13084
rect 11192 13028 11196 13084
rect 11132 13024 11196 13028
rect 17079 13084 17143 13088
rect 17079 13028 17083 13084
rect 17083 13028 17139 13084
rect 17139 13028 17143 13084
rect 17079 13024 17143 13028
rect 17159 13084 17223 13088
rect 17159 13028 17163 13084
rect 17163 13028 17219 13084
rect 17219 13028 17223 13084
rect 17159 13024 17223 13028
rect 17239 13084 17303 13088
rect 17239 13028 17243 13084
rect 17243 13028 17299 13084
rect 17299 13028 17303 13084
rect 17239 13024 17303 13028
rect 17319 13084 17383 13088
rect 17319 13028 17323 13084
rect 17323 13028 17379 13084
rect 17379 13028 17383 13084
rect 17319 13024 17383 13028
rect 23266 13084 23330 13088
rect 23266 13028 23270 13084
rect 23270 13028 23326 13084
rect 23326 13028 23330 13084
rect 23266 13024 23330 13028
rect 23346 13084 23410 13088
rect 23346 13028 23350 13084
rect 23350 13028 23406 13084
rect 23406 13028 23410 13084
rect 23346 13024 23410 13028
rect 23426 13084 23490 13088
rect 23426 13028 23430 13084
rect 23430 13028 23486 13084
rect 23486 13028 23490 13084
rect 23426 13024 23490 13028
rect 23506 13084 23570 13088
rect 23506 13028 23510 13084
rect 23510 13028 23566 13084
rect 23566 13028 23570 13084
rect 23506 13024 23570 13028
rect 4045 12540 4109 12544
rect 4045 12484 4049 12540
rect 4049 12484 4105 12540
rect 4105 12484 4109 12540
rect 4045 12480 4109 12484
rect 4125 12540 4189 12544
rect 4125 12484 4129 12540
rect 4129 12484 4185 12540
rect 4185 12484 4189 12540
rect 4125 12480 4189 12484
rect 4205 12540 4269 12544
rect 4205 12484 4209 12540
rect 4209 12484 4265 12540
rect 4265 12484 4269 12540
rect 4205 12480 4269 12484
rect 4285 12540 4349 12544
rect 4285 12484 4289 12540
rect 4289 12484 4345 12540
rect 4345 12484 4349 12540
rect 4285 12480 4349 12484
rect 10232 12540 10296 12544
rect 10232 12484 10236 12540
rect 10236 12484 10292 12540
rect 10292 12484 10296 12540
rect 10232 12480 10296 12484
rect 10312 12540 10376 12544
rect 10312 12484 10316 12540
rect 10316 12484 10372 12540
rect 10372 12484 10376 12540
rect 10312 12480 10376 12484
rect 10392 12540 10456 12544
rect 10392 12484 10396 12540
rect 10396 12484 10452 12540
rect 10452 12484 10456 12540
rect 10392 12480 10456 12484
rect 10472 12540 10536 12544
rect 10472 12484 10476 12540
rect 10476 12484 10532 12540
rect 10532 12484 10536 12540
rect 10472 12480 10536 12484
rect 16419 12540 16483 12544
rect 16419 12484 16423 12540
rect 16423 12484 16479 12540
rect 16479 12484 16483 12540
rect 16419 12480 16483 12484
rect 16499 12540 16563 12544
rect 16499 12484 16503 12540
rect 16503 12484 16559 12540
rect 16559 12484 16563 12540
rect 16499 12480 16563 12484
rect 16579 12540 16643 12544
rect 16579 12484 16583 12540
rect 16583 12484 16639 12540
rect 16639 12484 16643 12540
rect 16579 12480 16643 12484
rect 16659 12540 16723 12544
rect 16659 12484 16663 12540
rect 16663 12484 16719 12540
rect 16719 12484 16723 12540
rect 16659 12480 16723 12484
rect 22606 12540 22670 12544
rect 22606 12484 22610 12540
rect 22610 12484 22666 12540
rect 22666 12484 22670 12540
rect 22606 12480 22670 12484
rect 22686 12540 22750 12544
rect 22686 12484 22690 12540
rect 22690 12484 22746 12540
rect 22746 12484 22750 12540
rect 22686 12480 22750 12484
rect 22766 12540 22830 12544
rect 22766 12484 22770 12540
rect 22770 12484 22826 12540
rect 22826 12484 22830 12540
rect 22766 12480 22830 12484
rect 22846 12540 22910 12544
rect 22846 12484 22850 12540
rect 22850 12484 22906 12540
rect 22906 12484 22910 12540
rect 22846 12480 22910 12484
rect 4705 11996 4769 12000
rect 4705 11940 4709 11996
rect 4709 11940 4765 11996
rect 4765 11940 4769 11996
rect 4705 11936 4769 11940
rect 4785 11996 4849 12000
rect 4785 11940 4789 11996
rect 4789 11940 4845 11996
rect 4845 11940 4849 11996
rect 4785 11936 4849 11940
rect 4865 11996 4929 12000
rect 4865 11940 4869 11996
rect 4869 11940 4925 11996
rect 4925 11940 4929 11996
rect 4865 11936 4929 11940
rect 4945 11996 5009 12000
rect 4945 11940 4949 11996
rect 4949 11940 5005 11996
rect 5005 11940 5009 11996
rect 4945 11936 5009 11940
rect 10892 11996 10956 12000
rect 10892 11940 10896 11996
rect 10896 11940 10952 11996
rect 10952 11940 10956 11996
rect 10892 11936 10956 11940
rect 10972 11996 11036 12000
rect 10972 11940 10976 11996
rect 10976 11940 11032 11996
rect 11032 11940 11036 11996
rect 10972 11936 11036 11940
rect 11052 11996 11116 12000
rect 11052 11940 11056 11996
rect 11056 11940 11112 11996
rect 11112 11940 11116 11996
rect 11052 11936 11116 11940
rect 11132 11996 11196 12000
rect 11132 11940 11136 11996
rect 11136 11940 11192 11996
rect 11192 11940 11196 11996
rect 11132 11936 11196 11940
rect 17079 11996 17143 12000
rect 17079 11940 17083 11996
rect 17083 11940 17139 11996
rect 17139 11940 17143 11996
rect 17079 11936 17143 11940
rect 17159 11996 17223 12000
rect 17159 11940 17163 11996
rect 17163 11940 17219 11996
rect 17219 11940 17223 11996
rect 17159 11936 17223 11940
rect 17239 11996 17303 12000
rect 17239 11940 17243 11996
rect 17243 11940 17299 11996
rect 17299 11940 17303 11996
rect 17239 11936 17303 11940
rect 17319 11996 17383 12000
rect 17319 11940 17323 11996
rect 17323 11940 17379 11996
rect 17379 11940 17383 11996
rect 17319 11936 17383 11940
rect 23266 11996 23330 12000
rect 23266 11940 23270 11996
rect 23270 11940 23326 11996
rect 23326 11940 23330 11996
rect 23266 11936 23330 11940
rect 23346 11996 23410 12000
rect 23346 11940 23350 11996
rect 23350 11940 23406 11996
rect 23406 11940 23410 11996
rect 23346 11936 23410 11940
rect 23426 11996 23490 12000
rect 23426 11940 23430 11996
rect 23430 11940 23486 11996
rect 23486 11940 23490 11996
rect 23426 11936 23490 11940
rect 23506 11996 23570 12000
rect 23506 11940 23510 11996
rect 23510 11940 23566 11996
rect 23566 11940 23570 11996
rect 23506 11936 23570 11940
rect 15332 11596 15396 11660
rect 4045 11452 4109 11456
rect 4045 11396 4049 11452
rect 4049 11396 4105 11452
rect 4105 11396 4109 11452
rect 4045 11392 4109 11396
rect 4125 11452 4189 11456
rect 4125 11396 4129 11452
rect 4129 11396 4185 11452
rect 4185 11396 4189 11452
rect 4125 11392 4189 11396
rect 4205 11452 4269 11456
rect 4205 11396 4209 11452
rect 4209 11396 4265 11452
rect 4265 11396 4269 11452
rect 4205 11392 4269 11396
rect 4285 11452 4349 11456
rect 4285 11396 4289 11452
rect 4289 11396 4345 11452
rect 4345 11396 4349 11452
rect 4285 11392 4349 11396
rect 10232 11452 10296 11456
rect 10232 11396 10236 11452
rect 10236 11396 10292 11452
rect 10292 11396 10296 11452
rect 10232 11392 10296 11396
rect 10312 11452 10376 11456
rect 10312 11396 10316 11452
rect 10316 11396 10372 11452
rect 10372 11396 10376 11452
rect 10312 11392 10376 11396
rect 10392 11452 10456 11456
rect 10392 11396 10396 11452
rect 10396 11396 10452 11452
rect 10452 11396 10456 11452
rect 10392 11392 10456 11396
rect 10472 11452 10536 11456
rect 10472 11396 10476 11452
rect 10476 11396 10532 11452
rect 10532 11396 10536 11452
rect 10472 11392 10536 11396
rect 16419 11452 16483 11456
rect 16419 11396 16423 11452
rect 16423 11396 16479 11452
rect 16479 11396 16483 11452
rect 16419 11392 16483 11396
rect 16499 11452 16563 11456
rect 16499 11396 16503 11452
rect 16503 11396 16559 11452
rect 16559 11396 16563 11452
rect 16499 11392 16563 11396
rect 16579 11452 16643 11456
rect 16579 11396 16583 11452
rect 16583 11396 16639 11452
rect 16639 11396 16643 11452
rect 16579 11392 16643 11396
rect 16659 11452 16723 11456
rect 16659 11396 16663 11452
rect 16663 11396 16719 11452
rect 16719 11396 16723 11452
rect 16659 11392 16723 11396
rect 22606 11452 22670 11456
rect 22606 11396 22610 11452
rect 22610 11396 22666 11452
rect 22666 11396 22670 11452
rect 22606 11392 22670 11396
rect 22686 11452 22750 11456
rect 22686 11396 22690 11452
rect 22690 11396 22746 11452
rect 22746 11396 22750 11452
rect 22686 11392 22750 11396
rect 22766 11452 22830 11456
rect 22766 11396 22770 11452
rect 22770 11396 22826 11452
rect 22826 11396 22830 11452
rect 22766 11392 22830 11396
rect 22846 11452 22910 11456
rect 22846 11396 22850 11452
rect 22850 11396 22906 11452
rect 22906 11396 22910 11452
rect 22846 11392 22910 11396
rect 4705 10908 4769 10912
rect 4705 10852 4709 10908
rect 4709 10852 4765 10908
rect 4765 10852 4769 10908
rect 4705 10848 4769 10852
rect 4785 10908 4849 10912
rect 4785 10852 4789 10908
rect 4789 10852 4845 10908
rect 4845 10852 4849 10908
rect 4785 10848 4849 10852
rect 4865 10908 4929 10912
rect 4865 10852 4869 10908
rect 4869 10852 4925 10908
rect 4925 10852 4929 10908
rect 4865 10848 4929 10852
rect 4945 10908 5009 10912
rect 4945 10852 4949 10908
rect 4949 10852 5005 10908
rect 5005 10852 5009 10908
rect 4945 10848 5009 10852
rect 10892 10908 10956 10912
rect 10892 10852 10896 10908
rect 10896 10852 10952 10908
rect 10952 10852 10956 10908
rect 10892 10848 10956 10852
rect 10972 10908 11036 10912
rect 10972 10852 10976 10908
rect 10976 10852 11032 10908
rect 11032 10852 11036 10908
rect 10972 10848 11036 10852
rect 11052 10908 11116 10912
rect 11052 10852 11056 10908
rect 11056 10852 11112 10908
rect 11112 10852 11116 10908
rect 11052 10848 11116 10852
rect 11132 10908 11196 10912
rect 11132 10852 11136 10908
rect 11136 10852 11192 10908
rect 11192 10852 11196 10908
rect 11132 10848 11196 10852
rect 17079 10908 17143 10912
rect 17079 10852 17083 10908
rect 17083 10852 17139 10908
rect 17139 10852 17143 10908
rect 17079 10848 17143 10852
rect 17159 10908 17223 10912
rect 17159 10852 17163 10908
rect 17163 10852 17219 10908
rect 17219 10852 17223 10908
rect 17159 10848 17223 10852
rect 17239 10908 17303 10912
rect 17239 10852 17243 10908
rect 17243 10852 17299 10908
rect 17299 10852 17303 10908
rect 17239 10848 17303 10852
rect 17319 10908 17383 10912
rect 17319 10852 17323 10908
rect 17323 10852 17379 10908
rect 17379 10852 17383 10908
rect 17319 10848 17383 10852
rect 23266 10908 23330 10912
rect 23266 10852 23270 10908
rect 23270 10852 23326 10908
rect 23326 10852 23330 10908
rect 23266 10848 23330 10852
rect 23346 10908 23410 10912
rect 23346 10852 23350 10908
rect 23350 10852 23406 10908
rect 23406 10852 23410 10908
rect 23346 10848 23410 10852
rect 23426 10908 23490 10912
rect 23426 10852 23430 10908
rect 23430 10852 23486 10908
rect 23486 10852 23490 10908
rect 23426 10848 23490 10852
rect 23506 10908 23570 10912
rect 23506 10852 23510 10908
rect 23510 10852 23566 10908
rect 23566 10852 23570 10908
rect 23506 10848 23570 10852
rect 4045 10364 4109 10368
rect 4045 10308 4049 10364
rect 4049 10308 4105 10364
rect 4105 10308 4109 10364
rect 4045 10304 4109 10308
rect 4125 10364 4189 10368
rect 4125 10308 4129 10364
rect 4129 10308 4185 10364
rect 4185 10308 4189 10364
rect 4125 10304 4189 10308
rect 4205 10364 4269 10368
rect 4205 10308 4209 10364
rect 4209 10308 4265 10364
rect 4265 10308 4269 10364
rect 4205 10304 4269 10308
rect 4285 10364 4349 10368
rect 4285 10308 4289 10364
rect 4289 10308 4345 10364
rect 4345 10308 4349 10364
rect 4285 10304 4349 10308
rect 10232 10364 10296 10368
rect 10232 10308 10236 10364
rect 10236 10308 10292 10364
rect 10292 10308 10296 10364
rect 10232 10304 10296 10308
rect 10312 10364 10376 10368
rect 10312 10308 10316 10364
rect 10316 10308 10372 10364
rect 10372 10308 10376 10364
rect 10312 10304 10376 10308
rect 10392 10364 10456 10368
rect 10392 10308 10396 10364
rect 10396 10308 10452 10364
rect 10452 10308 10456 10364
rect 10392 10304 10456 10308
rect 10472 10364 10536 10368
rect 10472 10308 10476 10364
rect 10476 10308 10532 10364
rect 10532 10308 10536 10364
rect 10472 10304 10536 10308
rect 16419 10364 16483 10368
rect 16419 10308 16423 10364
rect 16423 10308 16479 10364
rect 16479 10308 16483 10364
rect 16419 10304 16483 10308
rect 16499 10364 16563 10368
rect 16499 10308 16503 10364
rect 16503 10308 16559 10364
rect 16559 10308 16563 10364
rect 16499 10304 16563 10308
rect 16579 10364 16643 10368
rect 16579 10308 16583 10364
rect 16583 10308 16639 10364
rect 16639 10308 16643 10364
rect 16579 10304 16643 10308
rect 16659 10364 16723 10368
rect 16659 10308 16663 10364
rect 16663 10308 16719 10364
rect 16719 10308 16723 10364
rect 16659 10304 16723 10308
rect 22606 10364 22670 10368
rect 22606 10308 22610 10364
rect 22610 10308 22666 10364
rect 22666 10308 22670 10364
rect 22606 10304 22670 10308
rect 22686 10364 22750 10368
rect 22686 10308 22690 10364
rect 22690 10308 22746 10364
rect 22746 10308 22750 10364
rect 22686 10304 22750 10308
rect 22766 10364 22830 10368
rect 22766 10308 22770 10364
rect 22770 10308 22826 10364
rect 22826 10308 22830 10364
rect 22766 10304 22830 10308
rect 22846 10364 22910 10368
rect 22846 10308 22850 10364
rect 22850 10308 22906 10364
rect 22906 10308 22910 10364
rect 22846 10304 22910 10308
rect 4705 9820 4769 9824
rect 4705 9764 4709 9820
rect 4709 9764 4765 9820
rect 4765 9764 4769 9820
rect 4705 9760 4769 9764
rect 4785 9820 4849 9824
rect 4785 9764 4789 9820
rect 4789 9764 4845 9820
rect 4845 9764 4849 9820
rect 4785 9760 4849 9764
rect 4865 9820 4929 9824
rect 4865 9764 4869 9820
rect 4869 9764 4925 9820
rect 4925 9764 4929 9820
rect 4865 9760 4929 9764
rect 4945 9820 5009 9824
rect 4945 9764 4949 9820
rect 4949 9764 5005 9820
rect 5005 9764 5009 9820
rect 4945 9760 5009 9764
rect 10892 9820 10956 9824
rect 10892 9764 10896 9820
rect 10896 9764 10952 9820
rect 10952 9764 10956 9820
rect 10892 9760 10956 9764
rect 10972 9820 11036 9824
rect 10972 9764 10976 9820
rect 10976 9764 11032 9820
rect 11032 9764 11036 9820
rect 10972 9760 11036 9764
rect 11052 9820 11116 9824
rect 11052 9764 11056 9820
rect 11056 9764 11112 9820
rect 11112 9764 11116 9820
rect 11052 9760 11116 9764
rect 11132 9820 11196 9824
rect 11132 9764 11136 9820
rect 11136 9764 11192 9820
rect 11192 9764 11196 9820
rect 11132 9760 11196 9764
rect 17079 9820 17143 9824
rect 17079 9764 17083 9820
rect 17083 9764 17139 9820
rect 17139 9764 17143 9820
rect 17079 9760 17143 9764
rect 17159 9820 17223 9824
rect 17159 9764 17163 9820
rect 17163 9764 17219 9820
rect 17219 9764 17223 9820
rect 17159 9760 17223 9764
rect 17239 9820 17303 9824
rect 17239 9764 17243 9820
rect 17243 9764 17299 9820
rect 17299 9764 17303 9820
rect 17239 9760 17303 9764
rect 17319 9820 17383 9824
rect 17319 9764 17323 9820
rect 17323 9764 17379 9820
rect 17379 9764 17383 9820
rect 17319 9760 17383 9764
rect 23266 9820 23330 9824
rect 23266 9764 23270 9820
rect 23270 9764 23326 9820
rect 23326 9764 23330 9820
rect 23266 9760 23330 9764
rect 23346 9820 23410 9824
rect 23346 9764 23350 9820
rect 23350 9764 23406 9820
rect 23406 9764 23410 9820
rect 23346 9760 23410 9764
rect 23426 9820 23490 9824
rect 23426 9764 23430 9820
rect 23430 9764 23486 9820
rect 23486 9764 23490 9820
rect 23426 9760 23490 9764
rect 23506 9820 23570 9824
rect 23506 9764 23510 9820
rect 23510 9764 23566 9820
rect 23566 9764 23570 9820
rect 23506 9760 23570 9764
rect 4045 9276 4109 9280
rect 4045 9220 4049 9276
rect 4049 9220 4105 9276
rect 4105 9220 4109 9276
rect 4045 9216 4109 9220
rect 4125 9276 4189 9280
rect 4125 9220 4129 9276
rect 4129 9220 4185 9276
rect 4185 9220 4189 9276
rect 4125 9216 4189 9220
rect 4205 9276 4269 9280
rect 4205 9220 4209 9276
rect 4209 9220 4265 9276
rect 4265 9220 4269 9276
rect 4205 9216 4269 9220
rect 4285 9276 4349 9280
rect 4285 9220 4289 9276
rect 4289 9220 4345 9276
rect 4345 9220 4349 9276
rect 4285 9216 4349 9220
rect 10232 9276 10296 9280
rect 10232 9220 10236 9276
rect 10236 9220 10292 9276
rect 10292 9220 10296 9276
rect 10232 9216 10296 9220
rect 10312 9276 10376 9280
rect 10312 9220 10316 9276
rect 10316 9220 10372 9276
rect 10372 9220 10376 9276
rect 10312 9216 10376 9220
rect 10392 9276 10456 9280
rect 10392 9220 10396 9276
rect 10396 9220 10452 9276
rect 10452 9220 10456 9276
rect 10392 9216 10456 9220
rect 10472 9276 10536 9280
rect 10472 9220 10476 9276
rect 10476 9220 10532 9276
rect 10532 9220 10536 9276
rect 10472 9216 10536 9220
rect 16419 9276 16483 9280
rect 16419 9220 16423 9276
rect 16423 9220 16479 9276
rect 16479 9220 16483 9276
rect 16419 9216 16483 9220
rect 16499 9276 16563 9280
rect 16499 9220 16503 9276
rect 16503 9220 16559 9276
rect 16559 9220 16563 9276
rect 16499 9216 16563 9220
rect 16579 9276 16643 9280
rect 16579 9220 16583 9276
rect 16583 9220 16639 9276
rect 16639 9220 16643 9276
rect 16579 9216 16643 9220
rect 16659 9276 16723 9280
rect 16659 9220 16663 9276
rect 16663 9220 16719 9276
rect 16719 9220 16723 9276
rect 16659 9216 16723 9220
rect 22606 9276 22670 9280
rect 22606 9220 22610 9276
rect 22610 9220 22666 9276
rect 22666 9220 22670 9276
rect 22606 9216 22670 9220
rect 22686 9276 22750 9280
rect 22686 9220 22690 9276
rect 22690 9220 22746 9276
rect 22746 9220 22750 9276
rect 22686 9216 22750 9220
rect 22766 9276 22830 9280
rect 22766 9220 22770 9276
rect 22770 9220 22826 9276
rect 22826 9220 22830 9276
rect 22766 9216 22830 9220
rect 22846 9276 22910 9280
rect 22846 9220 22850 9276
rect 22850 9220 22906 9276
rect 22906 9220 22910 9276
rect 22846 9216 22910 9220
rect 4705 8732 4769 8736
rect 4705 8676 4709 8732
rect 4709 8676 4765 8732
rect 4765 8676 4769 8732
rect 4705 8672 4769 8676
rect 4785 8732 4849 8736
rect 4785 8676 4789 8732
rect 4789 8676 4845 8732
rect 4845 8676 4849 8732
rect 4785 8672 4849 8676
rect 4865 8732 4929 8736
rect 4865 8676 4869 8732
rect 4869 8676 4925 8732
rect 4925 8676 4929 8732
rect 4865 8672 4929 8676
rect 4945 8732 5009 8736
rect 4945 8676 4949 8732
rect 4949 8676 5005 8732
rect 5005 8676 5009 8732
rect 4945 8672 5009 8676
rect 10892 8732 10956 8736
rect 10892 8676 10896 8732
rect 10896 8676 10952 8732
rect 10952 8676 10956 8732
rect 10892 8672 10956 8676
rect 10972 8732 11036 8736
rect 10972 8676 10976 8732
rect 10976 8676 11032 8732
rect 11032 8676 11036 8732
rect 10972 8672 11036 8676
rect 11052 8732 11116 8736
rect 11052 8676 11056 8732
rect 11056 8676 11112 8732
rect 11112 8676 11116 8732
rect 11052 8672 11116 8676
rect 11132 8732 11196 8736
rect 11132 8676 11136 8732
rect 11136 8676 11192 8732
rect 11192 8676 11196 8732
rect 11132 8672 11196 8676
rect 17079 8732 17143 8736
rect 17079 8676 17083 8732
rect 17083 8676 17139 8732
rect 17139 8676 17143 8732
rect 17079 8672 17143 8676
rect 17159 8732 17223 8736
rect 17159 8676 17163 8732
rect 17163 8676 17219 8732
rect 17219 8676 17223 8732
rect 17159 8672 17223 8676
rect 17239 8732 17303 8736
rect 17239 8676 17243 8732
rect 17243 8676 17299 8732
rect 17299 8676 17303 8732
rect 17239 8672 17303 8676
rect 17319 8732 17383 8736
rect 17319 8676 17323 8732
rect 17323 8676 17379 8732
rect 17379 8676 17383 8732
rect 17319 8672 17383 8676
rect 23266 8732 23330 8736
rect 23266 8676 23270 8732
rect 23270 8676 23326 8732
rect 23326 8676 23330 8732
rect 23266 8672 23330 8676
rect 23346 8732 23410 8736
rect 23346 8676 23350 8732
rect 23350 8676 23406 8732
rect 23406 8676 23410 8732
rect 23346 8672 23410 8676
rect 23426 8732 23490 8736
rect 23426 8676 23430 8732
rect 23430 8676 23486 8732
rect 23486 8676 23490 8732
rect 23426 8672 23490 8676
rect 23506 8732 23570 8736
rect 23506 8676 23510 8732
rect 23510 8676 23566 8732
rect 23566 8676 23570 8732
rect 23506 8672 23570 8676
rect 4045 8188 4109 8192
rect 4045 8132 4049 8188
rect 4049 8132 4105 8188
rect 4105 8132 4109 8188
rect 4045 8128 4109 8132
rect 4125 8188 4189 8192
rect 4125 8132 4129 8188
rect 4129 8132 4185 8188
rect 4185 8132 4189 8188
rect 4125 8128 4189 8132
rect 4205 8188 4269 8192
rect 4205 8132 4209 8188
rect 4209 8132 4265 8188
rect 4265 8132 4269 8188
rect 4205 8128 4269 8132
rect 4285 8188 4349 8192
rect 4285 8132 4289 8188
rect 4289 8132 4345 8188
rect 4345 8132 4349 8188
rect 4285 8128 4349 8132
rect 10232 8188 10296 8192
rect 10232 8132 10236 8188
rect 10236 8132 10292 8188
rect 10292 8132 10296 8188
rect 10232 8128 10296 8132
rect 10312 8188 10376 8192
rect 10312 8132 10316 8188
rect 10316 8132 10372 8188
rect 10372 8132 10376 8188
rect 10312 8128 10376 8132
rect 10392 8188 10456 8192
rect 10392 8132 10396 8188
rect 10396 8132 10452 8188
rect 10452 8132 10456 8188
rect 10392 8128 10456 8132
rect 10472 8188 10536 8192
rect 10472 8132 10476 8188
rect 10476 8132 10532 8188
rect 10532 8132 10536 8188
rect 10472 8128 10536 8132
rect 16419 8188 16483 8192
rect 16419 8132 16423 8188
rect 16423 8132 16479 8188
rect 16479 8132 16483 8188
rect 16419 8128 16483 8132
rect 16499 8188 16563 8192
rect 16499 8132 16503 8188
rect 16503 8132 16559 8188
rect 16559 8132 16563 8188
rect 16499 8128 16563 8132
rect 16579 8188 16643 8192
rect 16579 8132 16583 8188
rect 16583 8132 16639 8188
rect 16639 8132 16643 8188
rect 16579 8128 16643 8132
rect 16659 8188 16723 8192
rect 16659 8132 16663 8188
rect 16663 8132 16719 8188
rect 16719 8132 16723 8188
rect 16659 8128 16723 8132
rect 22606 8188 22670 8192
rect 22606 8132 22610 8188
rect 22610 8132 22666 8188
rect 22666 8132 22670 8188
rect 22606 8128 22670 8132
rect 22686 8188 22750 8192
rect 22686 8132 22690 8188
rect 22690 8132 22746 8188
rect 22746 8132 22750 8188
rect 22686 8128 22750 8132
rect 22766 8188 22830 8192
rect 22766 8132 22770 8188
rect 22770 8132 22826 8188
rect 22826 8132 22830 8188
rect 22766 8128 22830 8132
rect 22846 8188 22910 8192
rect 22846 8132 22850 8188
rect 22850 8132 22906 8188
rect 22906 8132 22910 8188
rect 22846 8128 22910 8132
rect 4705 7644 4769 7648
rect 4705 7588 4709 7644
rect 4709 7588 4765 7644
rect 4765 7588 4769 7644
rect 4705 7584 4769 7588
rect 4785 7644 4849 7648
rect 4785 7588 4789 7644
rect 4789 7588 4845 7644
rect 4845 7588 4849 7644
rect 4785 7584 4849 7588
rect 4865 7644 4929 7648
rect 4865 7588 4869 7644
rect 4869 7588 4925 7644
rect 4925 7588 4929 7644
rect 4865 7584 4929 7588
rect 4945 7644 5009 7648
rect 4945 7588 4949 7644
rect 4949 7588 5005 7644
rect 5005 7588 5009 7644
rect 4945 7584 5009 7588
rect 10892 7644 10956 7648
rect 10892 7588 10896 7644
rect 10896 7588 10952 7644
rect 10952 7588 10956 7644
rect 10892 7584 10956 7588
rect 10972 7644 11036 7648
rect 10972 7588 10976 7644
rect 10976 7588 11032 7644
rect 11032 7588 11036 7644
rect 10972 7584 11036 7588
rect 11052 7644 11116 7648
rect 11052 7588 11056 7644
rect 11056 7588 11112 7644
rect 11112 7588 11116 7644
rect 11052 7584 11116 7588
rect 11132 7644 11196 7648
rect 11132 7588 11136 7644
rect 11136 7588 11192 7644
rect 11192 7588 11196 7644
rect 11132 7584 11196 7588
rect 17079 7644 17143 7648
rect 17079 7588 17083 7644
rect 17083 7588 17139 7644
rect 17139 7588 17143 7644
rect 17079 7584 17143 7588
rect 17159 7644 17223 7648
rect 17159 7588 17163 7644
rect 17163 7588 17219 7644
rect 17219 7588 17223 7644
rect 17159 7584 17223 7588
rect 17239 7644 17303 7648
rect 17239 7588 17243 7644
rect 17243 7588 17299 7644
rect 17299 7588 17303 7644
rect 17239 7584 17303 7588
rect 17319 7644 17383 7648
rect 17319 7588 17323 7644
rect 17323 7588 17379 7644
rect 17379 7588 17383 7644
rect 17319 7584 17383 7588
rect 23266 7644 23330 7648
rect 23266 7588 23270 7644
rect 23270 7588 23326 7644
rect 23326 7588 23330 7644
rect 23266 7584 23330 7588
rect 23346 7644 23410 7648
rect 23346 7588 23350 7644
rect 23350 7588 23406 7644
rect 23406 7588 23410 7644
rect 23346 7584 23410 7588
rect 23426 7644 23490 7648
rect 23426 7588 23430 7644
rect 23430 7588 23486 7644
rect 23486 7588 23490 7644
rect 23426 7584 23490 7588
rect 23506 7644 23570 7648
rect 23506 7588 23510 7644
rect 23510 7588 23566 7644
rect 23566 7588 23570 7644
rect 23506 7584 23570 7588
rect 4045 7100 4109 7104
rect 4045 7044 4049 7100
rect 4049 7044 4105 7100
rect 4105 7044 4109 7100
rect 4045 7040 4109 7044
rect 4125 7100 4189 7104
rect 4125 7044 4129 7100
rect 4129 7044 4185 7100
rect 4185 7044 4189 7100
rect 4125 7040 4189 7044
rect 4205 7100 4269 7104
rect 4205 7044 4209 7100
rect 4209 7044 4265 7100
rect 4265 7044 4269 7100
rect 4205 7040 4269 7044
rect 4285 7100 4349 7104
rect 4285 7044 4289 7100
rect 4289 7044 4345 7100
rect 4345 7044 4349 7100
rect 4285 7040 4349 7044
rect 10232 7100 10296 7104
rect 10232 7044 10236 7100
rect 10236 7044 10292 7100
rect 10292 7044 10296 7100
rect 10232 7040 10296 7044
rect 10312 7100 10376 7104
rect 10312 7044 10316 7100
rect 10316 7044 10372 7100
rect 10372 7044 10376 7100
rect 10312 7040 10376 7044
rect 10392 7100 10456 7104
rect 10392 7044 10396 7100
rect 10396 7044 10452 7100
rect 10452 7044 10456 7100
rect 10392 7040 10456 7044
rect 10472 7100 10536 7104
rect 10472 7044 10476 7100
rect 10476 7044 10532 7100
rect 10532 7044 10536 7100
rect 10472 7040 10536 7044
rect 16419 7100 16483 7104
rect 16419 7044 16423 7100
rect 16423 7044 16479 7100
rect 16479 7044 16483 7100
rect 16419 7040 16483 7044
rect 16499 7100 16563 7104
rect 16499 7044 16503 7100
rect 16503 7044 16559 7100
rect 16559 7044 16563 7100
rect 16499 7040 16563 7044
rect 16579 7100 16643 7104
rect 16579 7044 16583 7100
rect 16583 7044 16639 7100
rect 16639 7044 16643 7100
rect 16579 7040 16643 7044
rect 16659 7100 16723 7104
rect 16659 7044 16663 7100
rect 16663 7044 16719 7100
rect 16719 7044 16723 7100
rect 16659 7040 16723 7044
rect 22606 7100 22670 7104
rect 22606 7044 22610 7100
rect 22610 7044 22666 7100
rect 22666 7044 22670 7100
rect 22606 7040 22670 7044
rect 22686 7100 22750 7104
rect 22686 7044 22690 7100
rect 22690 7044 22746 7100
rect 22746 7044 22750 7100
rect 22686 7040 22750 7044
rect 22766 7100 22830 7104
rect 22766 7044 22770 7100
rect 22770 7044 22826 7100
rect 22826 7044 22830 7100
rect 22766 7040 22830 7044
rect 22846 7100 22910 7104
rect 22846 7044 22850 7100
rect 22850 7044 22906 7100
rect 22906 7044 22910 7100
rect 22846 7040 22910 7044
rect 4705 6556 4769 6560
rect 4705 6500 4709 6556
rect 4709 6500 4765 6556
rect 4765 6500 4769 6556
rect 4705 6496 4769 6500
rect 4785 6556 4849 6560
rect 4785 6500 4789 6556
rect 4789 6500 4845 6556
rect 4845 6500 4849 6556
rect 4785 6496 4849 6500
rect 4865 6556 4929 6560
rect 4865 6500 4869 6556
rect 4869 6500 4925 6556
rect 4925 6500 4929 6556
rect 4865 6496 4929 6500
rect 4945 6556 5009 6560
rect 4945 6500 4949 6556
rect 4949 6500 5005 6556
rect 5005 6500 5009 6556
rect 4945 6496 5009 6500
rect 10892 6556 10956 6560
rect 10892 6500 10896 6556
rect 10896 6500 10952 6556
rect 10952 6500 10956 6556
rect 10892 6496 10956 6500
rect 10972 6556 11036 6560
rect 10972 6500 10976 6556
rect 10976 6500 11032 6556
rect 11032 6500 11036 6556
rect 10972 6496 11036 6500
rect 11052 6556 11116 6560
rect 11052 6500 11056 6556
rect 11056 6500 11112 6556
rect 11112 6500 11116 6556
rect 11052 6496 11116 6500
rect 11132 6556 11196 6560
rect 11132 6500 11136 6556
rect 11136 6500 11192 6556
rect 11192 6500 11196 6556
rect 11132 6496 11196 6500
rect 17079 6556 17143 6560
rect 17079 6500 17083 6556
rect 17083 6500 17139 6556
rect 17139 6500 17143 6556
rect 17079 6496 17143 6500
rect 17159 6556 17223 6560
rect 17159 6500 17163 6556
rect 17163 6500 17219 6556
rect 17219 6500 17223 6556
rect 17159 6496 17223 6500
rect 17239 6556 17303 6560
rect 17239 6500 17243 6556
rect 17243 6500 17299 6556
rect 17299 6500 17303 6556
rect 17239 6496 17303 6500
rect 17319 6556 17383 6560
rect 17319 6500 17323 6556
rect 17323 6500 17379 6556
rect 17379 6500 17383 6556
rect 17319 6496 17383 6500
rect 23266 6556 23330 6560
rect 23266 6500 23270 6556
rect 23270 6500 23326 6556
rect 23326 6500 23330 6556
rect 23266 6496 23330 6500
rect 23346 6556 23410 6560
rect 23346 6500 23350 6556
rect 23350 6500 23406 6556
rect 23406 6500 23410 6556
rect 23346 6496 23410 6500
rect 23426 6556 23490 6560
rect 23426 6500 23430 6556
rect 23430 6500 23486 6556
rect 23486 6500 23490 6556
rect 23426 6496 23490 6500
rect 23506 6556 23570 6560
rect 23506 6500 23510 6556
rect 23510 6500 23566 6556
rect 23566 6500 23570 6556
rect 23506 6496 23570 6500
rect 4045 6012 4109 6016
rect 4045 5956 4049 6012
rect 4049 5956 4105 6012
rect 4105 5956 4109 6012
rect 4045 5952 4109 5956
rect 4125 6012 4189 6016
rect 4125 5956 4129 6012
rect 4129 5956 4185 6012
rect 4185 5956 4189 6012
rect 4125 5952 4189 5956
rect 4205 6012 4269 6016
rect 4205 5956 4209 6012
rect 4209 5956 4265 6012
rect 4265 5956 4269 6012
rect 4205 5952 4269 5956
rect 4285 6012 4349 6016
rect 4285 5956 4289 6012
rect 4289 5956 4345 6012
rect 4345 5956 4349 6012
rect 4285 5952 4349 5956
rect 10232 6012 10296 6016
rect 10232 5956 10236 6012
rect 10236 5956 10292 6012
rect 10292 5956 10296 6012
rect 10232 5952 10296 5956
rect 10312 6012 10376 6016
rect 10312 5956 10316 6012
rect 10316 5956 10372 6012
rect 10372 5956 10376 6012
rect 10312 5952 10376 5956
rect 10392 6012 10456 6016
rect 10392 5956 10396 6012
rect 10396 5956 10452 6012
rect 10452 5956 10456 6012
rect 10392 5952 10456 5956
rect 10472 6012 10536 6016
rect 10472 5956 10476 6012
rect 10476 5956 10532 6012
rect 10532 5956 10536 6012
rect 10472 5952 10536 5956
rect 16419 6012 16483 6016
rect 16419 5956 16423 6012
rect 16423 5956 16479 6012
rect 16479 5956 16483 6012
rect 16419 5952 16483 5956
rect 16499 6012 16563 6016
rect 16499 5956 16503 6012
rect 16503 5956 16559 6012
rect 16559 5956 16563 6012
rect 16499 5952 16563 5956
rect 16579 6012 16643 6016
rect 16579 5956 16583 6012
rect 16583 5956 16639 6012
rect 16639 5956 16643 6012
rect 16579 5952 16643 5956
rect 16659 6012 16723 6016
rect 16659 5956 16663 6012
rect 16663 5956 16719 6012
rect 16719 5956 16723 6012
rect 16659 5952 16723 5956
rect 22606 6012 22670 6016
rect 22606 5956 22610 6012
rect 22610 5956 22666 6012
rect 22666 5956 22670 6012
rect 22606 5952 22670 5956
rect 22686 6012 22750 6016
rect 22686 5956 22690 6012
rect 22690 5956 22746 6012
rect 22746 5956 22750 6012
rect 22686 5952 22750 5956
rect 22766 6012 22830 6016
rect 22766 5956 22770 6012
rect 22770 5956 22826 6012
rect 22826 5956 22830 6012
rect 22766 5952 22830 5956
rect 22846 6012 22910 6016
rect 22846 5956 22850 6012
rect 22850 5956 22906 6012
rect 22906 5956 22910 6012
rect 22846 5952 22910 5956
rect 4705 5468 4769 5472
rect 4705 5412 4709 5468
rect 4709 5412 4765 5468
rect 4765 5412 4769 5468
rect 4705 5408 4769 5412
rect 4785 5468 4849 5472
rect 4785 5412 4789 5468
rect 4789 5412 4845 5468
rect 4845 5412 4849 5468
rect 4785 5408 4849 5412
rect 4865 5468 4929 5472
rect 4865 5412 4869 5468
rect 4869 5412 4925 5468
rect 4925 5412 4929 5468
rect 4865 5408 4929 5412
rect 4945 5468 5009 5472
rect 4945 5412 4949 5468
rect 4949 5412 5005 5468
rect 5005 5412 5009 5468
rect 4945 5408 5009 5412
rect 10892 5468 10956 5472
rect 10892 5412 10896 5468
rect 10896 5412 10952 5468
rect 10952 5412 10956 5468
rect 10892 5408 10956 5412
rect 10972 5468 11036 5472
rect 10972 5412 10976 5468
rect 10976 5412 11032 5468
rect 11032 5412 11036 5468
rect 10972 5408 11036 5412
rect 11052 5468 11116 5472
rect 11052 5412 11056 5468
rect 11056 5412 11112 5468
rect 11112 5412 11116 5468
rect 11052 5408 11116 5412
rect 11132 5468 11196 5472
rect 11132 5412 11136 5468
rect 11136 5412 11192 5468
rect 11192 5412 11196 5468
rect 11132 5408 11196 5412
rect 17079 5468 17143 5472
rect 17079 5412 17083 5468
rect 17083 5412 17139 5468
rect 17139 5412 17143 5468
rect 17079 5408 17143 5412
rect 17159 5468 17223 5472
rect 17159 5412 17163 5468
rect 17163 5412 17219 5468
rect 17219 5412 17223 5468
rect 17159 5408 17223 5412
rect 17239 5468 17303 5472
rect 17239 5412 17243 5468
rect 17243 5412 17299 5468
rect 17299 5412 17303 5468
rect 17239 5408 17303 5412
rect 17319 5468 17383 5472
rect 17319 5412 17323 5468
rect 17323 5412 17379 5468
rect 17379 5412 17383 5468
rect 17319 5408 17383 5412
rect 23266 5468 23330 5472
rect 23266 5412 23270 5468
rect 23270 5412 23326 5468
rect 23326 5412 23330 5468
rect 23266 5408 23330 5412
rect 23346 5468 23410 5472
rect 23346 5412 23350 5468
rect 23350 5412 23406 5468
rect 23406 5412 23410 5468
rect 23346 5408 23410 5412
rect 23426 5468 23490 5472
rect 23426 5412 23430 5468
rect 23430 5412 23486 5468
rect 23486 5412 23490 5468
rect 23426 5408 23490 5412
rect 23506 5468 23570 5472
rect 23506 5412 23510 5468
rect 23510 5412 23566 5468
rect 23566 5412 23570 5468
rect 23506 5408 23570 5412
rect 4045 4924 4109 4928
rect 4045 4868 4049 4924
rect 4049 4868 4105 4924
rect 4105 4868 4109 4924
rect 4045 4864 4109 4868
rect 4125 4924 4189 4928
rect 4125 4868 4129 4924
rect 4129 4868 4185 4924
rect 4185 4868 4189 4924
rect 4125 4864 4189 4868
rect 4205 4924 4269 4928
rect 4205 4868 4209 4924
rect 4209 4868 4265 4924
rect 4265 4868 4269 4924
rect 4205 4864 4269 4868
rect 4285 4924 4349 4928
rect 4285 4868 4289 4924
rect 4289 4868 4345 4924
rect 4345 4868 4349 4924
rect 4285 4864 4349 4868
rect 10232 4924 10296 4928
rect 10232 4868 10236 4924
rect 10236 4868 10292 4924
rect 10292 4868 10296 4924
rect 10232 4864 10296 4868
rect 10312 4924 10376 4928
rect 10312 4868 10316 4924
rect 10316 4868 10372 4924
rect 10372 4868 10376 4924
rect 10312 4864 10376 4868
rect 10392 4924 10456 4928
rect 10392 4868 10396 4924
rect 10396 4868 10452 4924
rect 10452 4868 10456 4924
rect 10392 4864 10456 4868
rect 10472 4924 10536 4928
rect 10472 4868 10476 4924
rect 10476 4868 10532 4924
rect 10532 4868 10536 4924
rect 10472 4864 10536 4868
rect 16419 4924 16483 4928
rect 16419 4868 16423 4924
rect 16423 4868 16479 4924
rect 16479 4868 16483 4924
rect 16419 4864 16483 4868
rect 16499 4924 16563 4928
rect 16499 4868 16503 4924
rect 16503 4868 16559 4924
rect 16559 4868 16563 4924
rect 16499 4864 16563 4868
rect 16579 4924 16643 4928
rect 16579 4868 16583 4924
rect 16583 4868 16639 4924
rect 16639 4868 16643 4924
rect 16579 4864 16643 4868
rect 16659 4924 16723 4928
rect 16659 4868 16663 4924
rect 16663 4868 16719 4924
rect 16719 4868 16723 4924
rect 16659 4864 16723 4868
rect 22606 4924 22670 4928
rect 22606 4868 22610 4924
rect 22610 4868 22666 4924
rect 22666 4868 22670 4924
rect 22606 4864 22670 4868
rect 22686 4924 22750 4928
rect 22686 4868 22690 4924
rect 22690 4868 22746 4924
rect 22746 4868 22750 4924
rect 22686 4864 22750 4868
rect 22766 4924 22830 4928
rect 22766 4868 22770 4924
rect 22770 4868 22826 4924
rect 22826 4868 22830 4924
rect 22766 4864 22830 4868
rect 22846 4924 22910 4928
rect 22846 4868 22850 4924
rect 22850 4868 22906 4924
rect 22906 4868 22910 4924
rect 22846 4864 22910 4868
rect 4705 4380 4769 4384
rect 4705 4324 4709 4380
rect 4709 4324 4765 4380
rect 4765 4324 4769 4380
rect 4705 4320 4769 4324
rect 4785 4380 4849 4384
rect 4785 4324 4789 4380
rect 4789 4324 4845 4380
rect 4845 4324 4849 4380
rect 4785 4320 4849 4324
rect 4865 4380 4929 4384
rect 4865 4324 4869 4380
rect 4869 4324 4925 4380
rect 4925 4324 4929 4380
rect 4865 4320 4929 4324
rect 4945 4380 5009 4384
rect 4945 4324 4949 4380
rect 4949 4324 5005 4380
rect 5005 4324 5009 4380
rect 4945 4320 5009 4324
rect 10892 4380 10956 4384
rect 10892 4324 10896 4380
rect 10896 4324 10952 4380
rect 10952 4324 10956 4380
rect 10892 4320 10956 4324
rect 10972 4380 11036 4384
rect 10972 4324 10976 4380
rect 10976 4324 11032 4380
rect 11032 4324 11036 4380
rect 10972 4320 11036 4324
rect 11052 4380 11116 4384
rect 11052 4324 11056 4380
rect 11056 4324 11112 4380
rect 11112 4324 11116 4380
rect 11052 4320 11116 4324
rect 11132 4380 11196 4384
rect 11132 4324 11136 4380
rect 11136 4324 11192 4380
rect 11192 4324 11196 4380
rect 11132 4320 11196 4324
rect 17079 4380 17143 4384
rect 17079 4324 17083 4380
rect 17083 4324 17139 4380
rect 17139 4324 17143 4380
rect 17079 4320 17143 4324
rect 17159 4380 17223 4384
rect 17159 4324 17163 4380
rect 17163 4324 17219 4380
rect 17219 4324 17223 4380
rect 17159 4320 17223 4324
rect 17239 4380 17303 4384
rect 17239 4324 17243 4380
rect 17243 4324 17299 4380
rect 17299 4324 17303 4380
rect 17239 4320 17303 4324
rect 17319 4380 17383 4384
rect 17319 4324 17323 4380
rect 17323 4324 17379 4380
rect 17379 4324 17383 4380
rect 17319 4320 17383 4324
rect 23266 4380 23330 4384
rect 23266 4324 23270 4380
rect 23270 4324 23326 4380
rect 23326 4324 23330 4380
rect 23266 4320 23330 4324
rect 23346 4380 23410 4384
rect 23346 4324 23350 4380
rect 23350 4324 23406 4380
rect 23406 4324 23410 4380
rect 23346 4320 23410 4324
rect 23426 4380 23490 4384
rect 23426 4324 23430 4380
rect 23430 4324 23486 4380
rect 23486 4324 23490 4380
rect 23426 4320 23490 4324
rect 23506 4380 23570 4384
rect 23506 4324 23510 4380
rect 23510 4324 23566 4380
rect 23566 4324 23570 4380
rect 23506 4320 23570 4324
rect 4045 3836 4109 3840
rect 4045 3780 4049 3836
rect 4049 3780 4105 3836
rect 4105 3780 4109 3836
rect 4045 3776 4109 3780
rect 4125 3836 4189 3840
rect 4125 3780 4129 3836
rect 4129 3780 4185 3836
rect 4185 3780 4189 3836
rect 4125 3776 4189 3780
rect 4205 3836 4269 3840
rect 4205 3780 4209 3836
rect 4209 3780 4265 3836
rect 4265 3780 4269 3836
rect 4205 3776 4269 3780
rect 4285 3836 4349 3840
rect 4285 3780 4289 3836
rect 4289 3780 4345 3836
rect 4345 3780 4349 3836
rect 4285 3776 4349 3780
rect 10232 3836 10296 3840
rect 10232 3780 10236 3836
rect 10236 3780 10292 3836
rect 10292 3780 10296 3836
rect 10232 3776 10296 3780
rect 10312 3836 10376 3840
rect 10312 3780 10316 3836
rect 10316 3780 10372 3836
rect 10372 3780 10376 3836
rect 10312 3776 10376 3780
rect 10392 3836 10456 3840
rect 10392 3780 10396 3836
rect 10396 3780 10452 3836
rect 10452 3780 10456 3836
rect 10392 3776 10456 3780
rect 10472 3836 10536 3840
rect 10472 3780 10476 3836
rect 10476 3780 10532 3836
rect 10532 3780 10536 3836
rect 10472 3776 10536 3780
rect 16419 3836 16483 3840
rect 16419 3780 16423 3836
rect 16423 3780 16479 3836
rect 16479 3780 16483 3836
rect 16419 3776 16483 3780
rect 16499 3836 16563 3840
rect 16499 3780 16503 3836
rect 16503 3780 16559 3836
rect 16559 3780 16563 3836
rect 16499 3776 16563 3780
rect 16579 3836 16643 3840
rect 16579 3780 16583 3836
rect 16583 3780 16639 3836
rect 16639 3780 16643 3836
rect 16579 3776 16643 3780
rect 16659 3836 16723 3840
rect 16659 3780 16663 3836
rect 16663 3780 16719 3836
rect 16719 3780 16723 3836
rect 16659 3776 16723 3780
rect 22606 3836 22670 3840
rect 22606 3780 22610 3836
rect 22610 3780 22666 3836
rect 22666 3780 22670 3836
rect 22606 3776 22670 3780
rect 22686 3836 22750 3840
rect 22686 3780 22690 3836
rect 22690 3780 22746 3836
rect 22746 3780 22750 3836
rect 22686 3776 22750 3780
rect 22766 3836 22830 3840
rect 22766 3780 22770 3836
rect 22770 3780 22826 3836
rect 22826 3780 22830 3836
rect 22766 3776 22830 3780
rect 22846 3836 22910 3840
rect 22846 3780 22850 3836
rect 22850 3780 22906 3836
rect 22906 3780 22910 3836
rect 22846 3776 22910 3780
rect 4705 3292 4769 3296
rect 4705 3236 4709 3292
rect 4709 3236 4765 3292
rect 4765 3236 4769 3292
rect 4705 3232 4769 3236
rect 4785 3292 4849 3296
rect 4785 3236 4789 3292
rect 4789 3236 4845 3292
rect 4845 3236 4849 3292
rect 4785 3232 4849 3236
rect 4865 3292 4929 3296
rect 4865 3236 4869 3292
rect 4869 3236 4925 3292
rect 4925 3236 4929 3292
rect 4865 3232 4929 3236
rect 4945 3292 5009 3296
rect 4945 3236 4949 3292
rect 4949 3236 5005 3292
rect 5005 3236 5009 3292
rect 4945 3232 5009 3236
rect 10892 3292 10956 3296
rect 10892 3236 10896 3292
rect 10896 3236 10952 3292
rect 10952 3236 10956 3292
rect 10892 3232 10956 3236
rect 10972 3292 11036 3296
rect 10972 3236 10976 3292
rect 10976 3236 11032 3292
rect 11032 3236 11036 3292
rect 10972 3232 11036 3236
rect 11052 3292 11116 3296
rect 11052 3236 11056 3292
rect 11056 3236 11112 3292
rect 11112 3236 11116 3292
rect 11052 3232 11116 3236
rect 11132 3292 11196 3296
rect 11132 3236 11136 3292
rect 11136 3236 11192 3292
rect 11192 3236 11196 3292
rect 11132 3232 11196 3236
rect 17079 3292 17143 3296
rect 17079 3236 17083 3292
rect 17083 3236 17139 3292
rect 17139 3236 17143 3292
rect 17079 3232 17143 3236
rect 17159 3292 17223 3296
rect 17159 3236 17163 3292
rect 17163 3236 17219 3292
rect 17219 3236 17223 3292
rect 17159 3232 17223 3236
rect 17239 3292 17303 3296
rect 17239 3236 17243 3292
rect 17243 3236 17299 3292
rect 17299 3236 17303 3292
rect 17239 3232 17303 3236
rect 17319 3292 17383 3296
rect 17319 3236 17323 3292
rect 17323 3236 17379 3292
rect 17379 3236 17383 3292
rect 17319 3232 17383 3236
rect 23266 3292 23330 3296
rect 23266 3236 23270 3292
rect 23270 3236 23326 3292
rect 23326 3236 23330 3292
rect 23266 3232 23330 3236
rect 23346 3292 23410 3296
rect 23346 3236 23350 3292
rect 23350 3236 23406 3292
rect 23406 3236 23410 3292
rect 23346 3232 23410 3236
rect 23426 3292 23490 3296
rect 23426 3236 23430 3292
rect 23430 3236 23486 3292
rect 23486 3236 23490 3292
rect 23426 3232 23490 3236
rect 23506 3292 23570 3296
rect 23506 3236 23510 3292
rect 23510 3236 23566 3292
rect 23566 3236 23570 3292
rect 23506 3232 23570 3236
rect 4045 2748 4109 2752
rect 4045 2692 4049 2748
rect 4049 2692 4105 2748
rect 4105 2692 4109 2748
rect 4045 2688 4109 2692
rect 4125 2748 4189 2752
rect 4125 2692 4129 2748
rect 4129 2692 4185 2748
rect 4185 2692 4189 2748
rect 4125 2688 4189 2692
rect 4205 2748 4269 2752
rect 4205 2692 4209 2748
rect 4209 2692 4265 2748
rect 4265 2692 4269 2748
rect 4205 2688 4269 2692
rect 4285 2748 4349 2752
rect 4285 2692 4289 2748
rect 4289 2692 4345 2748
rect 4345 2692 4349 2748
rect 4285 2688 4349 2692
rect 10232 2748 10296 2752
rect 10232 2692 10236 2748
rect 10236 2692 10292 2748
rect 10292 2692 10296 2748
rect 10232 2688 10296 2692
rect 10312 2748 10376 2752
rect 10312 2692 10316 2748
rect 10316 2692 10372 2748
rect 10372 2692 10376 2748
rect 10312 2688 10376 2692
rect 10392 2748 10456 2752
rect 10392 2692 10396 2748
rect 10396 2692 10452 2748
rect 10452 2692 10456 2748
rect 10392 2688 10456 2692
rect 10472 2748 10536 2752
rect 10472 2692 10476 2748
rect 10476 2692 10532 2748
rect 10532 2692 10536 2748
rect 10472 2688 10536 2692
rect 16419 2748 16483 2752
rect 16419 2692 16423 2748
rect 16423 2692 16479 2748
rect 16479 2692 16483 2748
rect 16419 2688 16483 2692
rect 16499 2748 16563 2752
rect 16499 2692 16503 2748
rect 16503 2692 16559 2748
rect 16559 2692 16563 2748
rect 16499 2688 16563 2692
rect 16579 2748 16643 2752
rect 16579 2692 16583 2748
rect 16583 2692 16639 2748
rect 16639 2692 16643 2748
rect 16579 2688 16643 2692
rect 16659 2748 16723 2752
rect 16659 2692 16663 2748
rect 16663 2692 16719 2748
rect 16719 2692 16723 2748
rect 16659 2688 16723 2692
rect 22606 2748 22670 2752
rect 22606 2692 22610 2748
rect 22610 2692 22666 2748
rect 22666 2692 22670 2748
rect 22606 2688 22670 2692
rect 22686 2748 22750 2752
rect 22686 2692 22690 2748
rect 22690 2692 22746 2748
rect 22746 2692 22750 2748
rect 22686 2688 22750 2692
rect 22766 2748 22830 2752
rect 22766 2692 22770 2748
rect 22770 2692 22826 2748
rect 22826 2692 22830 2748
rect 22766 2688 22830 2692
rect 22846 2748 22910 2752
rect 22846 2692 22850 2748
rect 22850 2692 22906 2748
rect 22906 2692 22910 2748
rect 22846 2688 22910 2692
rect 15332 2620 15396 2684
rect 4705 2204 4769 2208
rect 4705 2148 4709 2204
rect 4709 2148 4765 2204
rect 4765 2148 4769 2204
rect 4705 2144 4769 2148
rect 4785 2204 4849 2208
rect 4785 2148 4789 2204
rect 4789 2148 4845 2204
rect 4845 2148 4849 2204
rect 4785 2144 4849 2148
rect 4865 2204 4929 2208
rect 4865 2148 4869 2204
rect 4869 2148 4925 2204
rect 4925 2148 4929 2204
rect 4865 2144 4929 2148
rect 4945 2204 5009 2208
rect 4945 2148 4949 2204
rect 4949 2148 5005 2204
rect 5005 2148 5009 2204
rect 4945 2144 5009 2148
rect 10892 2204 10956 2208
rect 10892 2148 10896 2204
rect 10896 2148 10952 2204
rect 10952 2148 10956 2204
rect 10892 2144 10956 2148
rect 10972 2204 11036 2208
rect 10972 2148 10976 2204
rect 10976 2148 11032 2204
rect 11032 2148 11036 2204
rect 10972 2144 11036 2148
rect 11052 2204 11116 2208
rect 11052 2148 11056 2204
rect 11056 2148 11112 2204
rect 11112 2148 11116 2204
rect 11052 2144 11116 2148
rect 11132 2204 11196 2208
rect 11132 2148 11136 2204
rect 11136 2148 11192 2204
rect 11192 2148 11196 2204
rect 11132 2144 11196 2148
rect 17079 2204 17143 2208
rect 17079 2148 17083 2204
rect 17083 2148 17139 2204
rect 17139 2148 17143 2204
rect 17079 2144 17143 2148
rect 17159 2204 17223 2208
rect 17159 2148 17163 2204
rect 17163 2148 17219 2204
rect 17219 2148 17223 2204
rect 17159 2144 17223 2148
rect 17239 2204 17303 2208
rect 17239 2148 17243 2204
rect 17243 2148 17299 2204
rect 17299 2148 17303 2204
rect 17239 2144 17303 2148
rect 17319 2204 17383 2208
rect 17319 2148 17323 2204
rect 17323 2148 17379 2204
rect 17379 2148 17383 2204
rect 17319 2144 17383 2148
rect 23266 2204 23330 2208
rect 23266 2148 23270 2204
rect 23270 2148 23326 2204
rect 23326 2148 23330 2204
rect 23266 2144 23330 2148
rect 23346 2204 23410 2208
rect 23346 2148 23350 2204
rect 23350 2148 23406 2204
rect 23406 2148 23410 2204
rect 23346 2144 23410 2148
rect 23426 2204 23490 2208
rect 23426 2148 23430 2204
rect 23430 2148 23486 2204
rect 23486 2148 23490 2204
rect 23426 2144 23490 2148
rect 23506 2204 23570 2208
rect 23506 2148 23510 2204
rect 23510 2148 23566 2204
rect 23566 2148 23570 2204
rect 23506 2144 23570 2148
<< metal4 >>
rect 4037 26688 4357 26704
rect 4037 26624 4045 26688
rect 4109 26624 4125 26688
rect 4189 26624 4205 26688
rect 4269 26624 4285 26688
rect 4349 26624 4357 26688
rect 4037 25600 4357 26624
rect 4037 25536 4045 25600
rect 4109 25536 4125 25600
rect 4189 25536 4205 25600
rect 4269 25536 4285 25600
rect 4349 25536 4357 25600
rect 4037 24512 4357 25536
rect 4037 24448 4045 24512
rect 4109 24448 4125 24512
rect 4189 24448 4205 24512
rect 4269 24448 4285 24512
rect 4349 24448 4357 24512
rect 4037 23714 4357 24448
rect 4037 23478 4079 23714
rect 4315 23478 4357 23714
rect 4037 23424 4357 23478
rect 4037 23360 4045 23424
rect 4109 23360 4125 23424
rect 4189 23360 4205 23424
rect 4269 23360 4285 23424
rect 4349 23360 4357 23424
rect 4037 22336 4357 23360
rect 4037 22272 4045 22336
rect 4109 22272 4125 22336
rect 4189 22272 4205 22336
rect 4269 22272 4285 22336
rect 4349 22272 4357 22336
rect 4037 21248 4357 22272
rect 4037 21184 4045 21248
rect 4109 21184 4125 21248
rect 4189 21184 4205 21248
rect 4269 21184 4285 21248
rect 4349 21184 4357 21248
rect 4037 20160 4357 21184
rect 4037 20096 4045 20160
rect 4109 20096 4125 20160
rect 4189 20096 4205 20160
rect 4269 20096 4285 20160
rect 4349 20096 4357 20160
rect 4037 19072 4357 20096
rect 4037 19008 4045 19072
rect 4109 19008 4125 19072
rect 4189 19008 4205 19072
rect 4269 19008 4285 19072
rect 4349 19008 4357 19072
rect 4037 17984 4357 19008
rect 4037 17920 4045 17984
rect 4109 17920 4125 17984
rect 4189 17920 4205 17984
rect 4269 17920 4285 17984
rect 4349 17920 4357 17984
rect 4037 17594 4357 17920
rect 4037 17358 4079 17594
rect 4315 17358 4357 17594
rect 4037 16896 4357 17358
rect 4037 16832 4045 16896
rect 4109 16832 4125 16896
rect 4189 16832 4205 16896
rect 4269 16832 4285 16896
rect 4349 16832 4357 16896
rect 4037 15808 4357 16832
rect 4037 15744 4045 15808
rect 4109 15744 4125 15808
rect 4189 15744 4205 15808
rect 4269 15744 4285 15808
rect 4349 15744 4357 15808
rect 4037 14720 4357 15744
rect 4037 14656 4045 14720
rect 4109 14656 4125 14720
rect 4189 14656 4205 14720
rect 4269 14656 4285 14720
rect 4349 14656 4357 14720
rect 4037 13632 4357 14656
rect 4037 13568 4045 13632
rect 4109 13568 4125 13632
rect 4189 13568 4205 13632
rect 4269 13568 4285 13632
rect 4349 13568 4357 13632
rect 4037 12544 4357 13568
rect 4037 12480 4045 12544
rect 4109 12480 4125 12544
rect 4189 12480 4205 12544
rect 4269 12480 4285 12544
rect 4349 12480 4357 12544
rect 4037 11474 4357 12480
rect 4037 11456 4079 11474
rect 4315 11456 4357 11474
rect 4037 11392 4045 11456
rect 4349 11392 4357 11456
rect 4037 11238 4079 11392
rect 4315 11238 4357 11392
rect 4037 10368 4357 11238
rect 4037 10304 4045 10368
rect 4109 10304 4125 10368
rect 4189 10304 4205 10368
rect 4269 10304 4285 10368
rect 4349 10304 4357 10368
rect 4037 9280 4357 10304
rect 4037 9216 4045 9280
rect 4109 9216 4125 9280
rect 4189 9216 4205 9280
rect 4269 9216 4285 9280
rect 4349 9216 4357 9280
rect 4037 8192 4357 9216
rect 4037 8128 4045 8192
rect 4109 8128 4125 8192
rect 4189 8128 4205 8192
rect 4269 8128 4285 8192
rect 4349 8128 4357 8192
rect 4037 7104 4357 8128
rect 4037 7040 4045 7104
rect 4109 7040 4125 7104
rect 4189 7040 4205 7104
rect 4269 7040 4285 7104
rect 4349 7040 4357 7104
rect 4037 6016 4357 7040
rect 4037 5952 4045 6016
rect 4109 5952 4125 6016
rect 4189 5952 4205 6016
rect 4269 5952 4285 6016
rect 4349 5952 4357 6016
rect 4037 5354 4357 5952
rect 4037 5118 4079 5354
rect 4315 5118 4357 5354
rect 4037 4928 4357 5118
rect 4037 4864 4045 4928
rect 4109 4864 4125 4928
rect 4189 4864 4205 4928
rect 4269 4864 4285 4928
rect 4349 4864 4357 4928
rect 4037 3840 4357 4864
rect 4037 3776 4045 3840
rect 4109 3776 4125 3840
rect 4189 3776 4205 3840
rect 4269 3776 4285 3840
rect 4349 3776 4357 3840
rect 4037 2752 4357 3776
rect 4037 2688 4045 2752
rect 4109 2688 4125 2752
rect 4189 2688 4205 2752
rect 4269 2688 4285 2752
rect 4349 2688 4357 2752
rect 4037 2128 4357 2688
rect 4697 26144 5017 26704
rect 4697 26080 4705 26144
rect 4769 26080 4785 26144
rect 4849 26080 4865 26144
rect 4929 26080 4945 26144
rect 5009 26080 5017 26144
rect 4697 25056 5017 26080
rect 4697 24992 4705 25056
rect 4769 24992 4785 25056
rect 4849 24992 4865 25056
rect 4929 24992 4945 25056
rect 5009 24992 5017 25056
rect 4697 24374 5017 24992
rect 10224 26688 10544 26704
rect 10224 26624 10232 26688
rect 10296 26624 10312 26688
rect 10376 26624 10392 26688
rect 10456 26624 10472 26688
rect 10536 26624 10544 26688
rect 10224 25600 10544 26624
rect 10224 25536 10232 25600
rect 10296 25536 10312 25600
rect 10376 25536 10392 25600
rect 10456 25536 10472 25600
rect 10536 25536 10544 25600
rect 9811 24716 9877 24717
rect 9811 24652 9812 24716
rect 9876 24652 9877 24716
rect 9811 24651 9877 24652
rect 4697 24138 4739 24374
rect 4975 24138 5017 24374
rect 4697 23968 5017 24138
rect 4697 23904 4705 23968
rect 4769 23904 4785 23968
rect 4849 23904 4865 23968
rect 4929 23904 4945 23968
rect 5009 23904 5017 23968
rect 4697 22880 5017 23904
rect 4697 22816 4705 22880
rect 4769 22816 4785 22880
rect 4849 22816 4865 22880
rect 4929 22816 4945 22880
rect 5009 22816 5017 22880
rect 4697 21792 5017 22816
rect 9814 22813 9874 24651
rect 10224 24512 10544 25536
rect 10224 24448 10232 24512
rect 10296 24448 10312 24512
rect 10376 24448 10392 24512
rect 10456 24448 10472 24512
rect 10536 24448 10544 24512
rect 10224 23714 10544 24448
rect 10224 23478 10266 23714
rect 10502 23478 10544 23714
rect 10224 23424 10544 23478
rect 10224 23360 10232 23424
rect 10296 23360 10312 23424
rect 10376 23360 10392 23424
rect 10456 23360 10472 23424
rect 10536 23360 10544 23424
rect 9811 22812 9877 22813
rect 9811 22748 9812 22812
rect 9876 22748 9877 22812
rect 9811 22747 9877 22748
rect 4697 21728 4705 21792
rect 4769 21728 4785 21792
rect 4849 21728 4865 21792
rect 4929 21728 4945 21792
rect 5009 21728 5017 21792
rect 4697 20704 5017 21728
rect 10224 22336 10544 23360
rect 10224 22272 10232 22336
rect 10296 22272 10312 22336
rect 10376 22272 10392 22336
rect 10456 22272 10472 22336
rect 10536 22272 10544 22336
rect 10224 21248 10544 22272
rect 10224 21184 10232 21248
rect 10296 21184 10312 21248
rect 10376 21184 10392 21248
rect 10456 21184 10472 21248
rect 10536 21184 10544 21248
rect 7787 20772 7853 20773
rect 7787 20708 7788 20772
rect 7852 20708 7853 20772
rect 7787 20707 7853 20708
rect 4697 20640 4705 20704
rect 4769 20640 4785 20704
rect 4849 20640 4865 20704
rect 4929 20640 4945 20704
rect 5009 20640 5017 20704
rect 4697 19616 5017 20640
rect 4697 19552 4705 19616
rect 4769 19552 4785 19616
rect 4849 19552 4865 19616
rect 4929 19552 4945 19616
rect 5009 19552 5017 19616
rect 4697 18528 5017 19552
rect 4697 18464 4705 18528
rect 4769 18464 4785 18528
rect 4849 18464 4865 18528
rect 4929 18464 4945 18528
rect 5009 18464 5017 18528
rect 4697 18254 5017 18464
rect 4697 18018 4739 18254
rect 4975 18018 5017 18254
rect 4697 17440 5017 18018
rect 7790 17917 7850 20707
rect 10224 20160 10544 21184
rect 10224 20096 10232 20160
rect 10296 20096 10312 20160
rect 10376 20096 10392 20160
rect 10456 20096 10472 20160
rect 10536 20096 10544 20160
rect 10224 19072 10544 20096
rect 10224 19008 10232 19072
rect 10296 19008 10312 19072
rect 10376 19008 10392 19072
rect 10456 19008 10472 19072
rect 10536 19008 10544 19072
rect 10224 17984 10544 19008
rect 10224 17920 10232 17984
rect 10296 17920 10312 17984
rect 10376 17920 10392 17984
rect 10456 17920 10472 17984
rect 10536 17920 10544 17984
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 4697 17376 4705 17440
rect 4769 17376 4785 17440
rect 4849 17376 4865 17440
rect 4929 17376 4945 17440
rect 5009 17376 5017 17440
rect 4697 16352 5017 17376
rect 4697 16288 4705 16352
rect 4769 16288 4785 16352
rect 4849 16288 4865 16352
rect 4929 16288 4945 16352
rect 5009 16288 5017 16352
rect 4697 15264 5017 16288
rect 4697 15200 4705 15264
rect 4769 15200 4785 15264
rect 4849 15200 4865 15264
rect 4929 15200 4945 15264
rect 5009 15200 5017 15264
rect 4697 14176 5017 15200
rect 4697 14112 4705 14176
rect 4769 14112 4785 14176
rect 4849 14112 4865 14176
rect 4929 14112 4945 14176
rect 5009 14112 5017 14176
rect 4697 13088 5017 14112
rect 4697 13024 4705 13088
rect 4769 13024 4785 13088
rect 4849 13024 4865 13088
rect 4929 13024 4945 13088
rect 5009 13024 5017 13088
rect 4697 12134 5017 13024
rect 4697 12000 4739 12134
rect 4975 12000 5017 12134
rect 4697 11936 4705 12000
rect 5009 11936 5017 12000
rect 4697 11898 4739 11936
rect 4975 11898 5017 11936
rect 4697 10912 5017 11898
rect 4697 10848 4705 10912
rect 4769 10848 4785 10912
rect 4849 10848 4865 10912
rect 4929 10848 4945 10912
rect 5009 10848 5017 10912
rect 4697 9824 5017 10848
rect 4697 9760 4705 9824
rect 4769 9760 4785 9824
rect 4849 9760 4865 9824
rect 4929 9760 4945 9824
rect 5009 9760 5017 9824
rect 4697 8736 5017 9760
rect 4697 8672 4705 8736
rect 4769 8672 4785 8736
rect 4849 8672 4865 8736
rect 4929 8672 4945 8736
rect 5009 8672 5017 8736
rect 4697 7648 5017 8672
rect 4697 7584 4705 7648
rect 4769 7584 4785 7648
rect 4849 7584 4865 7648
rect 4929 7584 4945 7648
rect 5009 7584 5017 7648
rect 4697 6560 5017 7584
rect 4697 6496 4705 6560
rect 4769 6496 4785 6560
rect 4849 6496 4865 6560
rect 4929 6496 4945 6560
rect 5009 6496 5017 6560
rect 4697 6014 5017 6496
rect 4697 5778 4739 6014
rect 4975 5778 5017 6014
rect 4697 5472 5017 5778
rect 4697 5408 4705 5472
rect 4769 5408 4785 5472
rect 4849 5408 4865 5472
rect 4929 5408 4945 5472
rect 5009 5408 5017 5472
rect 4697 4384 5017 5408
rect 4697 4320 4705 4384
rect 4769 4320 4785 4384
rect 4849 4320 4865 4384
rect 4929 4320 4945 4384
rect 5009 4320 5017 4384
rect 4697 3296 5017 4320
rect 4697 3232 4705 3296
rect 4769 3232 4785 3296
rect 4849 3232 4865 3296
rect 4929 3232 4945 3296
rect 5009 3232 5017 3296
rect 4697 2208 5017 3232
rect 4697 2144 4705 2208
rect 4769 2144 4785 2208
rect 4849 2144 4865 2208
rect 4929 2144 4945 2208
rect 5009 2144 5017 2208
rect 4697 2128 5017 2144
rect 10224 17594 10544 17920
rect 10224 17358 10266 17594
rect 10502 17358 10544 17594
rect 10224 16896 10544 17358
rect 10224 16832 10232 16896
rect 10296 16832 10312 16896
rect 10376 16832 10392 16896
rect 10456 16832 10472 16896
rect 10536 16832 10544 16896
rect 10224 15808 10544 16832
rect 10224 15744 10232 15808
rect 10296 15744 10312 15808
rect 10376 15744 10392 15808
rect 10456 15744 10472 15808
rect 10536 15744 10544 15808
rect 10224 14720 10544 15744
rect 10224 14656 10232 14720
rect 10296 14656 10312 14720
rect 10376 14656 10392 14720
rect 10456 14656 10472 14720
rect 10536 14656 10544 14720
rect 10224 13632 10544 14656
rect 10224 13568 10232 13632
rect 10296 13568 10312 13632
rect 10376 13568 10392 13632
rect 10456 13568 10472 13632
rect 10536 13568 10544 13632
rect 10224 12544 10544 13568
rect 10224 12480 10232 12544
rect 10296 12480 10312 12544
rect 10376 12480 10392 12544
rect 10456 12480 10472 12544
rect 10536 12480 10544 12544
rect 10224 11474 10544 12480
rect 10224 11456 10266 11474
rect 10502 11456 10544 11474
rect 10224 11392 10232 11456
rect 10536 11392 10544 11456
rect 10224 11238 10266 11392
rect 10502 11238 10544 11392
rect 10224 10368 10544 11238
rect 10224 10304 10232 10368
rect 10296 10304 10312 10368
rect 10376 10304 10392 10368
rect 10456 10304 10472 10368
rect 10536 10304 10544 10368
rect 10224 9280 10544 10304
rect 10224 9216 10232 9280
rect 10296 9216 10312 9280
rect 10376 9216 10392 9280
rect 10456 9216 10472 9280
rect 10536 9216 10544 9280
rect 10224 8192 10544 9216
rect 10224 8128 10232 8192
rect 10296 8128 10312 8192
rect 10376 8128 10392 8192
rect 10456 8128 10472 8192
rect 10536 8128 10544 8192
rect 10224 7104 10544 8128
rect 10224 7040 10232 7104
rect 10296 7040 10312 7104
rect 10376 7040 10392 7104
rect 10456 7040 10472 7104
rect 10536 7040 10544 7104
rect 10224 6016 10544 7040
rect 10224 5952 10232 6016
rect 10296 5952 10312 6016
rect 10376 5952 10392 6016
rect 10456 5952 10472 6016
rect 10536 5952 10544 6016
rect 10224 5354 10544 5952
rect 10224 5118 10266 5354
rect 10502 5118 10544 5354
rect 10224 4928 10544 5118
rect 10224 4864 10232 4928
rect 10296 4864 10312 4928
rect 10376 4864 10392 4928
rect 10456 4864 10472 4928
rect 10536 4864 10544 4928
rect 10224 3840 10544 4864
rect 10224 3776 10232 3840
rect 10296 3776 10312 3840
rect 10376 3776 10392 3840
rect 10456 3776 10472 3840
rect 10536 3776 10544 3840
rect 10224 2752 10544 3776
rect 10224 2688 10232 2752
rect 10296 2688 10312 2752
rect 10376 2688 10392 2752
rect 10456 2688 10472 2752
rect 10536 2688 10544 2752
rect 10224 2128 10544 2688
rect 10884 26144 11204 26704
rect 10884 26080 10892 26144
rect 10956 26080 10972 26144
rect 11036 26080 11052 26144
rect 11116 26080 11132 26144
rect 11196 26080 11204 26144
rect 10884 25056 11204 26080
rect 10884 24992 10892 25056
rect 10956 24992 10972 25056
rect 11036 24992 11052 25056
rect 11116 24992 11132 25056
rect 11196 24992 11204 25056
rect 10884 24374 11204 24992
rect 10884 24138 10926 24374
rect 11162 24138 11204 24374
rect 10884 23968 11204 24138
rect 10884 23904 10892 23968
rect 10956 23904 10972 23968
rect 11036 23904 11052 23968
rect 11116 23904 11132 23968
rect 11196 23904 11204 23968
rect 10884 22880 11204 23904
rect 10884 22816 10892 22880
rect 10956 22816 10972 22880
rect 11036 22816 11052 22880
rect 11116 22816 11132 22880
rect 11196 22816 11204 22880
rect 10884 21792 11204 22816
rect 10884 21728 10892 21792
rect 10956 21728 10972 21792
rect 11036 21728 11052 21792
rect 11116 21728 11132 21792
rect 11196 21728 11204 21792
rect 10884 20704 11204 21728
rect 10884 20640 10892 20704
rect 10956 20640 10972 20704
rect 11036 20640 11052 20704
rect 11116 20640 11132 20704
rect 11196 20640 11204 20704
rect 10884 19616 11204 20640
rect 10884 19552 10892 19616
rect 10956 19552 10972 19616
rect 11036 19552 11052 19616
rect 11116 19552 11132 19616
rect 11196 19552 11204 19616
rect 10884 18528 11204 19552
rect 10884 18464 10892 18528
rect 10956 18464 10972 18528
rect 11036 18464 11052 18528
rect 11116 18464 11132 18528
rect 11196 18464 11204 18528
rect 10884 18254 11204 18464
rect 10884 18018 10926 18254
rect 11162 18018 11204 18254
rect 10884 17440 11204 18018
rect 10884 17376 10892 17440
rect 10956 17376 10972 17440
rect 11036 17376 11052 17440
rect 11116 17376 11132 17440
rect 11196 17376 11204 17440
rect 10884 16352 11204 17376
rect 10884 16288 10892 16352
rect 10956 16288 10972 16352
rect 11036 16288 11052 16352
rect 11116 16288 11132 16352
rect 11196 16288 11204 16352
rect 10884 15264 11204 16288
rect 10884 15200 10892 15264
rect 10956 15200 10972 15264
rect 11036 15200 11052 15264
rect 11116 15200 11132 15264
rect 11196 15200 11204 15264
rect 10884 14176 11204 15200
rect 10884 14112 10892 14176
rect 10956 14112 10972 14176
rect 11036 14112 11052 14176
rect 11116 14112 11132 14176
rect 11196 14112 11204 14176
rect 10884 13088 11204 14112
rect 10884 13024 10892 13088
rect 10956 13024 10972 13088
rect 11036 13024 11052 13088
rect 11116 13024 11132 13088
rect 11196 13024 11204 13088
rect 10884 12134 11204 13024
rect 10884 12000 10926 12134
rect 11162 12000 11204 12134
rect 10884 11936 10892 12000
rect 11196 11936 11204 12000
rect 10884 11898 10926 11936
rect 11162 11898 11204 11936
rect 10884 10912 11204 11898
rect 16411 26688 16731 26704
rect 16411 26624 16419 26688
rect 16483 26624 16499 26688
rect 16563 26624 16579 26688
rect 16643 26624 16659 26688
rect 16723 26624 16731 26688
rect 16411 25600 16731 26624
rect 16411 25536 16419 25600
rect 16483 25536 16499 25600
rect 16563 25536 16579 25600
rect 16643 25536 16659 25600
rect 16723 25536 16731 25600
rect 16411 24512 16731 25536
rect 16411 24448 16419 24512
rect 16483 24448 16499 24512
rect 16563 24448 16579 24512
rect 16643 24448 16659 24512
rect 16723 24448 16731 24512
rect 16411 23714 16731 24448
rect 16411 23478 16453 23714
rect 16689 23478 16731 23714
rect 16411 23424 16731 23478
rect 16411 23360 16419 23424
rect 16483 23360 16499 23424
rect 16563 23360 16579 23424
rect 16643 23360 16659 23424
rect 16723 23360 16731 23424
rect 16411 22336 16731 23360
rect 16411 22272 16419 22336
rect 16483 22272 16499 22336
rect 16563 22272 16579 22336
rect 16643 22272 16659 22336
rect 16723 22272 16731 22336
rect 16411 21248 16731 22272
rect 16411 21184 16419 21248
rect 16483 21184 16499 21248
rect 16563 21184 16579 21248
rect 16643 21184 16659 21248
rect 16723 21184 16731 21248
rect 16411 20160 16731 21184
rect 16411 20096 16419 20160
rect 16483 20096 16499 20160
rect 16563 20096 16579 20160
rect 16643 20096 16659 20160
rect 16723 20096 16731 20160
rect 16411 19072 16731 20096
rect 16411 19008 16419 19072
rect 16483 19008 16499 19072
rect 16563 19008 16579 19072
rect 16643 19008 16659 19072
rect 16723 19008 16731 19072
rect 16411 17984 16731 19008
rect 16411 17920 16419 17984
rect 16483 17920 16499 17984
rect 16563 17920 16579 17984
rect 16643 17920 16659 17984
rect 16723 17920 16731 17984
rect 16411 17594 16731 17920
rect 16411 17358 16453 17594
rect 16689 17358 16731 17594
rect 16411 16896 16731 17358
rect 16411 16832 16419 16896
rect 16483 16832 16499 16896
rect 16563 16832 16579 16896
rect 16643 16832 16659 16896
rect 16723 16832 16731 16896
rect 16411 15808 16731 16832
rect 16411 15744 16419 15808
rect 16483 15744 16499 15808
rect 16563 15744 16579 15808
rect 16643 15744 16659 15808
rect 16723 15744 16731 15808
rect 16411 14720 16731 15744
rect 16411 14656 16419 14720
rect 16483 14656 16499 14720
rect 16563 14656 16579 14720
rect 16643 14656 16659 14720
rect 16723 14656 16731 14720
rect 16411 13632 16731 14656
rect 16411 13568 16419 13632
rect 16483 13568 16499 13632
rect 16563 13568 16579 13632
rect 16643 13568 16659 13632
rect 16723 13568 16731 13632
rect 16411 12544 16731 13568
rect 16411 12480 16419 12544
rect 16483 12480 16499 12544
rect 16563 12480 16579 12544
rect 16643 12480 16659 12544
rect 16723 12480 16731 12544
rect 15331 11660 15397 11661
rect 15331 11596 15332 11660
rect 15396 11596 15397 11660
rect 15331 11595 15397 11596
rect 10884 10848 10892 10912
rect 10956 10848 10972 10912
rect 11036 10848 11052 10912
rect 11116 10848 11132 10912
rect 11196 10848 11204 10912
rect 10884 9824 11204 10848
rect 10884 9760 10892 9824
rect 10956 9760 10972 9824
rect 11036 9760 11052 9824
rect 11116 9760 11132 9824
rect 11196 9760 11204 9824
rect 10884 8736 11204 9760
rect 10884 8672 10892 8736
rect 10956 8672 10972 8736
rect 11036 8672 11052 8736
rect 11116 8672 11132 8736
rect 11196 8672 11204 8736
rect 10884 7648 11204 8672
rect 10884 7584 10892 7648
rect 10956 7584 10972 7648
rect 11036 7584 11052 7648
rect 11116 7584 11132 7648
rect 11196 7584 11204 7648
rect 10884 6560 11204 7584
rect 10884 6496 10892 6560
rect 10956 6496 10972 6560
rect 11036 6496 11052 6560
rect 11116 6496 11132 6560
rect 11196 6496 11204 6560
rect 10884 6014 11204 6496
rect 10884 5778 10926 6014
rect 11162 5778 11204 6014
rect 10884 5472 11204 5778
rect 10884 5408 10892 5472
rect 10956 5408 10972 5472
rect 11036 5408 11052 5472
rect 11116 5408 11132 5472
rect 11196 5408 11204 5472
rect 10884 4384 11204 5408
rect 10884 4320 10892 4384
rect 10956 4320 10972 4384
rect 11036 4320 11052 4384
rect 11116 4320 11132 4384
rect 11196 4320 11204 4384
rect 10884 3296 11204 4320
rect 10884 3232 10892 3296
rect 10956 3232 10972 3296
rect 11036 3232 11052 3296
rect 11116 3232 11132 3296
rect 11196 3232 11204 3296
rect 10884 2208 11204 3232
rect 15334 2685 15394 11595
rect 16411 11474 16731 12480
rect 16411 11456 16453 11474
rect 16689 11456 16731 11474
rect 16411 11392 16419 11456
rect 16723 11392 16731 11456
rect 16411 11238 16453 11392
rect 16689 11238 16731 11392
rect 16411 10368 16731 11238
rect 16411 10304 16419 10368
rect 16483 10304 16499 10368
rect 16563 10304 16579 10368
rect 16643 10304 16659 10368
rect 16723 10304 16731 10368
rect 16411 9280 16731 10304
rect 16411 9216 16419 9280
rect 16483 9216 16499 9280
rect 16563 9216 16579 9280
rect 16643 9216 16659 9280
rect 16723 9216 16731 9280
rect 16411 8192 16731 9216
rect 16411 8128 16419 8192
rect 16483 8128 16499 8192
rect 16563 8128 16579 8192
rect 16643 8128 16659 8192
rect 16723 8128 16731 8192
rect 16411 7104 16731 8128
rect 16411 7040 16419 7104
rect 16483 7040 16499 7104
rect 16563 7040 16579 7104
rect 16643 7040 16659 7104
rect 16723 7040 16731 7104
rect 16411 6016 16731 7040
rect 16411 5952 16419 6016
rect 16483 5952 16499 6016
rect 16563 5952 16579 6016
rect 16643 5952 16659 6016
rect 16723 5952 16731 6016
rect 16411 5354 16731 5952
rect 16411 5118 16453 5354
rect 16689 5118 16731 5354
rect 16411 4928 16731 5118
rect 16411 4864 16419 4928
rect 16483 4864 16499 4928
rect 16563 4864 16579 4928
rect 16643 4864 16659 4928
rect 16723 4864 16731 4928
rect 16411 3840 16731 4864
rect 16411 3776 16419 3840
rect 16483 3776 16499 3840
rect 16563 3776 16579 3840
rect 16643 3776 16659 3840
rect 16723 3776 16731 3840
rect 16411 2752 16731 3776
rect 16411 2688 16419 2752
rect 16483 2688 16499 2752
rect 16563 2688 16579 2752
rect 16643 2688 16659 2752
rect 16723 2688 16731 2752
rect 15331 2684 15397 2685
rect 15331 2620 15332 2684
rect 15396 2620 15397 2684
rect 15331 2619 15397 2620
rect 10884 2144 10892 2208
rect 10956 2144 10972 2208
rect 11036 2144 11052 2208
rect 11116 2144 11132 2208
rect 11196 2144 11204 2208
rect 10884 2128 11204 2144
rect 16411 2128 16731 2688
rect 17071 26144 17391 26704
rect 17071 26080 17079 26144
rect 17143 26080 17159 26144
rect 17223 26080 17239 26144
rect 17303 26080 17319 26144
rect 17383 26080 17391 26144
rect 17071 25056 17391 26080
rect 17071 24992 17079 25056
rect 17143 24992 17159 25056
rect 17223 24992 17239 25056
rect 17303 24992 17319 25056
rect 17383 24992 17391 25056
rect 17071 24374 17391 24992
rect 17071 24138 17113 24374
rect 17349 24138 17391 24374
rect 17071 23968 17391 24138
rect 17071 23904 17079 23968
rect 17143 23904 17159 23968
rect 17223 23904 17239 23968
rect 17303 23904 17319 23968
rect 17383 23904 17391 23968
rect 17071 22880 17391 23904
rect 17071 22816 17079 22880
rect 17143 22816 17159 22880
rect 17223 22816 17239 22880
rect 17303 22816 17319 22880
rect 17383 22816 17391 22880
rect 17071 21792 17391 22816
rect 17071 21728 17079 21792
rect 17143 21728 17159 21792
rect 17223 21728 17239 21792
rect 17303 21728 17319 21792
rect 17383 21728 17391 21792
rect 17071 20704 17391 21728
rect 17071 20640 17079 20704
rect 17143 20640 17159 20704
rect 17223 20640 17239 20704
rect 17303 20640 17319 20704
rect 17383 20640 17391 20704
rect 17071 19616 17391 20640
rect 17071 19552 17079 19616
rect 17143 19552 17159 19616
rect 17223 19552 17239 19616
rect 17303 19552 17319 19616
rect 17383 19552 17391 19616
rect 17071 18528 17391 19552
rect 17071 18464 17079 18528
rect 17143 18464 17159 18528
rect 17223 18464 17239 18528
rect 17303 18464 17319 18528
rect 17383 18464 17391 18528
rect 17071 18254 17391 18464
rect 17071 18018 17113 18254
rect 17349 18018 17391 18254
rect 17071 17440 17391 18018
rect 17071 17376 17079 17440
rect 17143 17376 17159 17440
rect 17223 17376 17239 17440
rect 17303 17376 17319 17440
rect 17383 17376 17391 17440
rect 17071 16352 17391 17376
rect 17071 16288 17079 16352
rect 17143 16288 17159 16352
rect 17223 16288 17239 16352
rect 17303 16288 17319 16352
rect 17383 16288 17391 16352
rect 17071 15264 17391 16288
rect 17071 15200 17079 15264
rect 17143 15200 17159 15264
rect 17223 15200 17239 15264
rect 17303 15200 17319 15264
rect 17383 15200 17391 15264
rect 17071 14176 17391 15200
rect 17071 14112 17079 14176
rect 17143 14112 17159 14176
rect 17223 14112 17239 14176
rect 17303 14112 17319 14176
rect 17383 14112 17391 14176
rect 17071 13088 17391 14112
rect 17071 13024 17079 13088
rect 17143 13024 17159 13088
rect 17223 13024 17239 13088
rect 17303 13024 17319 13088
rect 17383 13024 17391 13088
rect 17071 12134 17391 13024
rect 17071 12000 17113 12134
rect 17349 12000 17391 12134
rect 17071 11936 17079 12000
rect 17383 11936 17391 12000
rect 17071 11898 17113 11936
rect 17349 11898 17391 11936
rect 17071 10912 17391 11898
rect 17071 10848 17079 10912
rect 17143 10848 17159 10912
rect 17223 10848 17239 10912
rect 17303 10848 17319 10912
rect 17383 10848 17391 10912
rect 17071 9824 17391 10848
rect 17071 9760 17079 9824
rect 17143 9760 17159 9824
rect 17223 9760 17239 9824
rect 17303 9760 17319 9824
rect 17383 9760 17391 9824
rect 17071 8736 17391 9760
rect 17071 8672 17079 8736
rect 17143 8672 17159 8736
rect 17223 8672 17239 8736
rect 17303 8672 17319 8736
rect 17383 8672 17391 8736
rect 17071 7648 17391 8672
rect 17071 7584 17079 7648
rect 17143 7584 17159 7648
rect 17223 7584 17239 7648
rect 17303 7584 17319 7648
rect 17383 7584 17391 7648
rect 17071 6560 17391 7584
rect 17071 6496 17079 6560
rect 17143 6496 17159 6560
rect 17223 6496 17239 6560
rect 17303 6496 17319 6560
rect 17383 6496 17391 6560
rect 17071 6014 17391 6496
rect 17071 5778 17113 6014
rect 17349 5778 17391 6014
rect 17071 5472 17391 5778
rect 17071 5408 17079 5472
rect 17143 5408 17159 5472
rect 17223 5408 17239 5472
rect 17303 5408 17319 5472
rect 17383 5408 17391 5472
rect 17071 4384 17391 5408
rect 17071 4320 17079 4384
rect 17143 4320 17159 4384
rect 17223 4320 17239 4384
rect 17303 4320 17319 4384
rect 17383 4320 17391 4384
rect 17071 3296 17391 4320
rect 17071 3232 17079 3296
rect 17143 3232 17159 3296
rect 17223 3232 17239 3296
rect 17303 3232 17319 3296
rect 17383 3232 17391 3296
rect 17071 2208 17391 3232
rect 17071 2144 17079 2208
rect 17143 2144 17159 2208
rect 17223 2144 17239 2208
rect 17303 2144 17319 2208
rect 17383 2144 17391 2208
rect 17071 2128 17391 2144
rect 22598 26688 22918 26704
rect 22598 26624 22606 26688
rect 22670 26624 22686 26688
rect 22750 26624 22766 26688
rect 22830 26624 22846 26688
rect 22910 26624 22918 26688
rect 22598 25600 22918 26624
rect 22598 25536 22606 25600
rect 22670 25536 22686 25600
rect 22750 25536 22766 25600
rect 22830 25536 22846 25600
rect 22910 25536 22918 25600
rect 22598 24512 22918 25536
rect 22598 24448 22606 24512
rect 22670 24448 22686 24512
rect 22750 24448 22766 24512
rect 22830 24448 22846 24512
rect 22910 24448 22918 24512
rect 22598 23714 22918 24448
rect 22598 23478 22640 23714
rect 22876 23478 22918 23714
rect 22598 23424 22918 23478
rect 22598 23360 22606 23424
rect 22670 23360 22686 23424
rect 22750 23360 22766 23424
rect 22830 23360 22846 23424
rect 22910 23360 22918 23424
rect 22598 22336 22918 23360
rect 22598 22272 22606 22336
rect 22670 22272 22686 22336
rect 22750 22272 22766 22336
rect 22830 22272 22846 22336
rect 22910 22272 22918 22336
rect 22598 21248 22918 22272
rect 22598 21184 22606 21248
rect 22670 21184 22686 21248
rect 22750 21184 22766 21248
rect 22830 21184 22846 21248
rect 22910 21184 22918 21248
rect 22598 20160 22918 21184
rect 22598 20096 22606 20160
rect 22670 20096 22686 20160
rect 22750 20096 22766 20160
rect 22830 20096 22846 20160
rect 22910 20096 22918 20160
rect 22598 19072 22918 20096
rect 22598 19008 22606 19072
rect 22670 19008 22686 19072
rect 22750 19008 22766 19072
rect 22830 19008 22846 19072
rect 22910 19008 22918 19072
rect 22598 17984 22918 19008
rect 22598 17920 22606 17984
rect 22670 17920 22686 17984
rect 22750 17920 22766 17984
rect 22830 17920 22846 17984
rect 22910 17920 22918 17984
rect 22598 17594 22918 17920
rect 22598 17358 22640 17594
rect 22876 17358 22918 17594
rect 22598 16896 22918 17358
rect 22598 16832 22606 16896
rect 22670 16832 22686 16896
rect 22750 16832 22766 16896
rect 22830 16832 22846 16896
rect 22910 16832 22918 16896
rect 22598 15808 22918 16832
rect 22598 15744 22606 15808
rect 22670 15744 22686 15808
rect 22750 15744 22766 15808
rect 22830 15744 22846 15808
rect 22910 15744 22918 15808
rect 22598 14720 22918 15744
rect 22598 14656 22606 14720
rect 22670 14656 22686 14720
rect 22750 14656 22766 14720
rect 22830 14656 22846 14720
rect 22910 14656 22918 14720
rect 22598 13632 22918 14656
rect 22598 13568 22606 13632
rect 22670 13568 22686 13632
rect 22750 13568 22766 13632
rect 22830 13568 22846 13632
rect 22910 13568 22918 13632
rect 22598 12544 22918 13568
rect 22598 12480 22606 12544
rect 22670 12480 22686 12544
rect 22750 12480 22766 12544
rect 22830 12480 22846 12544
rect 22910 12480 22918 12544
rect 22598 11474 22918 12480
rect 22598 11456 22640 11474
rect 22876 11456 22918 11474
rect 22598 11392 22606 11456
rect 22910 11392 22918 11456
rect 22598 11238 22640 11392
rect 22876 11238 22918 11392
rect 22598 10368 22918 11238
rect 22598 10304 22606 10368
rect 22670 10304 22686 10368
rect 22750 10304 22766 10368
rect 22830 10304 22846 10368
rect 22910 10304 22918 10368
rect 22598 9280 22918 10304
rect 22598 9216 22606 9280
rect 22670 9216 22686 9280
rect 22750 9216 22766 9280
rect 22830 9216 22846 9280
rect 22910 9216 22918 9280
rect 22598 8192 22918 9216
rect 22598 8128 22606 8192
rect 22670 8128 22686 8192
rect 22750 8128 22766 8192
rect 22830 8128 22846 8192
rect 22910 8128 22918 8192
rect 22598 7104 22918 8128
rect 22598 7040 22606 7104
rect 22670 7040 22686 7104
rect 22750 7040 22766 7104
rect 22830 7040 22846 7104
rect 22910 7040 22918 7104
rect 22598 6016 22918 7040
rect 22598 5952 22606 6016
rect 22670 5952 22686 6016
rect 22750 5952 22766 6016
rect 22830 5952 22846 6016
rect 22910 5952 22918 6016
rect 22598 5354 22918 5952
rect 22598 5118 22640 5354
rect 22876 5118 22918 5354
rect 22598 4928 22918 5118
rect 22598 4864 22606 4928
rect 22670 4864 22686 4928
rect 22750 4864 22766 4928
rect 22830 4864 22846 4928
rect 22910 4864 22918 4928
rect 22598 3840 22918 4864
rect 22598 3776 22606 3840
rect 22670 3776 22686 3840
rect 22750 3776 22766 3840
rect 22830 3776 22846 3840
rect 22910 3776 22918 3840
rect 22598 2752 22918 3776
rect 22598 2688 22606 2752
rect 22670 2688 22686 2752
rect 22750 2688 22766 2752
rect 22830 2688 22846 2752
rect 22910 2688 22918 2752
rect 22598 2128 22918 2688
rect 23258 26144 23578 26704
rect 23258 26080 23266 26144
rect 23330 26080 23346 26144
rect 23410 26080 23426 26144
rect 23490 26080 23506 26144
rect 23570 26080 23578 26144
rect 23258 25056 23578 26080
rect 23258 24992 23266 25056
rect 23330 24992 23346 25056
rect 23410 24992 23426 25056
rect 23490 24992 23506 25056
rect 23570 24992 23578 25056
rect 23258 24374 23578 24992
rect 23258 24138 23300 24374
rect 23536 24138 23578 24374
rect 23258 23968 23578 24138
rect 23258 23904 23266 23968
rect 23330 23904 23346 23968
rect 23410 23904 23426 23968
rect 23490 23904 23506 23968
rect 23570 23904 23578 23968
rect 23258 22880 23578 23904
rect 23258 22816 23266 22880
rect 23330 22816 23346 22880
rect 23410 22816 23426 22880
rect 23490 22816 23506 22880
rect 23570 22816 23578 22880
rect 23258 21792 23578 22816
rect 23258 21728 23266 21792
rect 23330 21728 23346 21792
rect 23410 21728 23426 21792
rect 23490 21728 23506 21792
rect 23570 21728 23578 21792
rect 23258 20704 23578 21728
rect 23258 20640 23266 20704
rect 23330 20640 23346 20704
rect 23410 20640 23426 20704
rect 23490 20640 23506 20704
rect 23570 20640 23578 20704
rect 23258 19616 23578 20640
rect 23258 19552 23266 19616
rect 23330 19552 23346 19616
rect 23410 19552 23426 19616
rect 23490 19552 23506 19616
rect 23570 19552 23578 19616
rect 23258 18528 23578 19552
rect 23258 18464 23266 18528
rect 23330 18464 23346 18528
rect 23410 18464 23426 18528
rect 23490 18464 23506 18528
rect 23570 18464 23578 18528
rect 23258 18254 23578 18464
rect 23258 18018 23300 18254
rect 23536 18018 23578 18254
rect 23258 17440 23578 18018
rect 23258 17376 23266 17440
rect 23330 17376 23346 17440
rect 23410 17376 23426 17440
rect 23490 17376 23506 17440
rect 23570 17376 23578 17440
rect 23258 16352 23578 17376
rect 23258 16288 23266 16352
rect 23330 16288 23346 16352
rect 23410 16288 23426 16352
rect 23490 16288 23506 16352
rect 23570 16288 23578 16352
rect 23258 15264 23578 16288
rect 23258 15200 23266 15264
rect 23330 15200 23346 15264
rect 23410 15200 23426 15264
rect 23490 15200 23506 15264
rect 23570 15200 23578 15264
rect 23258 14176 23578 15200
rect 23258 14112 23266 14176
rect 23330 14112 23346 14176
rect 23410 14112 23426 14176
rect 23490 14112 23506 14176
rect 23570 14112 23578 14176
rect 23258 13088 23578 14112
rect 23258 13024 23266 13088
rect 23330 13024 23346 13088
rect 23410 13024 23426 13088
rect 23490 13024 23506 13088
rect 23570 13024 23578 13088
rect 23258 12134 23578 13024
rect 23258 12000 23300 12134
rect 23536 12000 23578 12134
rect 23258 11936 23266 12000
rect 23570 11936 23578 12000
rect 23258 11898 23300 11936
rect 23536 11898 23578 11936
rect 23258 10912 23578 11898
rect 23258 10848 23266 10912
rect 23330 10848 23346 10912
rect 23410 10848 23426 10912
rect 23490 10848 23506 10912
rect 23570 10848 23578 10912
rect 23258 9824 23578 10848
rect 23258 9760 23266 9824
rect 23330 9760 23346 9824
rect 23410 9760 23426 9824
rect 23490 9760 23506 9824
rect 23570 9760 23578 9824
rect 23258 8736 23578 9760
rect 23258 8672 23266 8736
rect 23330 8672 23346 8736
rect 23410 8672 23426 8736
rect 23490 8672 23506 8736
rect 23570 8672 23578 8736
rect 23258 7648 23578 8672
rect 23258 7584 23266 7648
rect 23330 7584 23346 7648
rect 23410 7584 23426 7648
rect 23490 7584 23506 7648
rect 23570 7584 23578 7648
rect 23258 6560 23578 7584
rect 23258 6496 23266 6560
rect 23330 6496 23346 6560
rect 23410 6496 23426 6560
rect 23490 6496 23506 6560
rect 23570 6496 23578 6560
rect 23258 6014 23578 6496
rect 23258 5778 23300 6014
rect 23536 5778 23578 6014
rect 23258 5472 23578 5778
rect 23258 5408 23266 5472
rect 23330 5408 23346 5472
rect 23410 5408 23426 5472
rect 23490 5408 23506 5472
rect 23570 5408 23578 5472
rect 23258 4384 23578 5408
rect 23258 4320 23266 4384
rect 23330 4320 23346 4384
rect 23410 4320 23426 4384
rect 23490 4320 23506 4384
rect 23570 4320 23578 4384
rect 23258 3296 23578 4320
rect 23258 3232 23266 3296
rect 23330 3232 23346 3296
rect 23410 3232 23426 3296
rect 23490 3232 23506 3296
rect 23570 3232 23578 3296
rect 23258 2208 23578 3232
rect 23258 2144 23266 2208
rect 23330 2144 23346 2208
rect 23410 2144 23426 2208
rect 23490 2144 23506 2208
rect 23570 2144 23578 2208
rect 23258 2128 23578 2144
<< via4 >>
rect 4079 23478 4315 23714
rect 4079 17358 4315 17594
rect 4079 11456 4315 11474
rect 4079 11392 4109 11456
rect 4109 11392 4125 11456
rect 4125 11392 4189 11456
rect 4189 11392 4205 11456
rect 4205 11392 4269 11456
rect 4269 11392 4285 11456
rect 4285 11392 4315 11456
rect 4079 11238 4315 11392
rect 4079 5118 4315 5354
rect 4739 24138 4975 24374
rect 10266 23478 10502 23714
rect 4739 18018 4975 18254
rect 4739 12000 4975 12134
rect 4739 11936 4769 12000
rect 4769 11936 4785 12000
rect 4785 11936 4849 12000
rect 4849 11936 4865 12000
rect 4865 11936 4929 12000
rect 4929 11936 4945 12000
rect 4945 11936 4975 12000
rect 4739 11898 4975 11936
rect 4739 5778 4975 6014
rect 10266 17358 10502 17594
rect 10266 11456 10502 11474
rect 10266 11392 10296 11456
rect 10296 11392 10312 11456
rect 10312 11392 10376 11456
rect 10376 11392 10392 11456
rect 10392 11392 10456 11456
rect 10456 11392 10472 11456
rect 10472 11392 10502 11456
rect 10266 11238 10502 11392
rect 10266 5118 10502 5354
rect 10926 24138 11162 24374
rect 10926 18018 11162 18254
rect 10926 12000 11162 12134
rect 10926 11936 10956 12000
rect 10956 11936 10972 12000
rect 10972 11936 11036 12000
rect 11036 11936 11052 12000
rect 11052 11936 11116 12000
rect 11116 11936 11132 12000
rect 11132 11936 11162 12000
rect 10926 11898 11162 11936
rect 16453 23478 16689 23714
rect 16453 17358 16689 17594
rect 10926 5778 11162 6014
rect 16453 11456 16689 11474
rect 16453 11392 16483 11456
rect 16483 11392 16499 11456
rect 16499 11392 16563 11456
rect 16563 11392 16579 11456
rect 16579 11392 16643 11456
rect 16643 11392 16659 11456
rect 16659 11392 16689 11456
rect 16453 11238 16689 11392
rect 16453 5118 16689 5354
rect 17113 24138 17349 24374
rect 17113 18018 17349 18254
rect 17113 12000 17349 12134
rect 17113 11936 17143 12000
rect 17143 11936 17159 12000
rect 17159 11936 17223 12000
rect 17223 11936 17239 12000
rect 17239 11936 17303 12000
rect 17303 11936 17319 12000
rect 17319 11936 17349 12000
rect 17113 11898 17349 11936
rect 17113 5778 17349 6014
rect 22640 23478 22876 23714
rect 22640 17358 22876 17594
rect 22640 11456 22876 11474
rect 22640 11392 22670 11456
rect 22670 11392 22686 11456
rect 22686 11392 22750 11456
rect 22750 11392 22766 11456
rect 22766 11392 22830 11456
rect 22830 11392 22846 11456
rect 22846 11392 22876 11456
rect 22640 11238 22876 11392
rect 22640 5118 22876 5354
rect 23300 24138 23536 24374
rect 23300 18018 23536 18254
rect 23300 12000 23536 12134
rect 23300 11936 23330 12000
rect 23330 11936 23346 12000
rect 23346 11936 23410 12000
rect 23410 11936 23426 12000
rect 23426 11936 23490 12000
rect 23490 11936 23506 12000
rect 23506 11936 23536 12000
rect 23300 11898 23536 11936
rect 23300 5778 23536 6014
<< metal5 >>
rect 1056 24374 25900 24416
rect 1056 24138 4739 24374
rect 4975 24138 10926 24374
rect 11162 24138 17113 24374
rect 17349 24138 23300 24374
rect 23536 24138 25900 24374
rect 1056 24096 25900 24138
rect 1056 23714 25900 23756
rect 1056 23478 4079 23714
rect 4315 23478 10266 23714
rect 10502 23478 16453 23714
rect 16689 23478 22640 23714
rect 22876 23478 25900 23714
rect 1056 23436 25900 23478
rect 1056 18254 25900 18296
rect 1056 18018 4739 18254
rect 4975 18018 10926 18254
rect 11162 18018 17113 18254
rect 17349 18018 23300 18254
rect 23536 18018 25900 18254
rect 1056 17976 25900 18018
rect 1056 17594 25900 17636
rect 1056 17358 4079 17594
rect 4315 17358 10266 17594
rect 10502 17358 16453 17594
rect 16689 17358 22640 17594
rect 22876 17358 25900 17594
rect 1056 17316 25900 17358
rect 1056 12134 25900 12176
rect 1056 11898 4739 12134
rect 4975 11898 10926 12134
rect 11162 11898 17113 12134
rect 17349 11898 23300 12134
rect 23536 11898 25900 12134
rect 1056 11856 25900 11898
rect 1056 11474 25900 11516
rect 1056 11238 4079 11474
rect 4315 11238 10266 11474
rect 10502 11238 16453 11474
rect 16689 11238 22640 11474
rect 22876 11238 25900 11474
rect 1056 11196 25900 11238
rect 1056 6014 25900 6056
rect 1056 5778 4739 6014
rect 4975 5778 10926 6014
rect 11162 5778 17113 6014
rect 17349 5778 23300 6014
rect 23536 5778 25900 6014
rect 1056 5736 25900 5778
rect 1056 5354 25900 5396
rect 1056 5118 4079 5354
rect 4315 5118 10266 5354
rect 10502 5118 16453 5354
rect 16689 5118 22640 5354
rect 22876 5118 25900 5354
rect 1056 5076 25900 5118
use sky130_fd_sc_hd__clkbuf_4  _0593_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0594_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0595_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1688980957
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0601_
timestamp 1688980957
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0604_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform 1 0 18216 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1688980957
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1688980957
transform 1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1688980957
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform 1 0 3128 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1688980957
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0625_
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform 1 0 6808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform 1 0 10580 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1688980957
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform 1 0 11960 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform 1 0 11960 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1688980957
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 1688980957
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1688980957
transform 1 0 21344 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0641_
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1688980957
transform 1 0 2392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0646_
timestamp 1688980957
transform 1 0 18032 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1688980957
transform 1 0 2944 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1688980957
transform 1 0 2392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0651_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0653_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1688980957
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0661_
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0662_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0664_
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0665_
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0666_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0667_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0668_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0669_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0670_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0672_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0673_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0675_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0676_
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0677_
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1688980957
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0679_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0680_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0681_
timestamp 1688980957
transform 1 0 8004 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_2  _0682_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0683_
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0685_
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0686_
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1688980957
transform 1 0 7544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0689_
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0690_
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0691_
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0692_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0693_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0694_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0695_
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0696_
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0697_
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0698_
timestamp 1688980957
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0699_
timestamp 1688980957
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0700_
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0701_
timestamp 1688980957
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0702_
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0704_
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0705_
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0707_
timestamp 1688980957
transform 1 0 19136 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0708_
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0709_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0710_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0711_
timestamp 1688980957
transform 1 0 7728 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0712_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o311ai_2  _0713_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0714_
timestamp 1688980957
transform 1 0 6532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0715_
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0716_
timestamp 1688980957
transform 1 0 6440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0717_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0718_
timestamp 1688980957
transform 1 0 4784 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0719_
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1688980957
transform 1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0721_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0722_
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0723_
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1688980957
transform 1 0 6992 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0725_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0727_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0728_
timestamp 1688980957
transform 1 0 5336 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0729_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0730_
timestamp 1688980957
transform 1 0 6440 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0731_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0732_
timestamp 1688980957
transform 1 0 14260 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0733_
timestamp 1688980957
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0734_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0735_
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _0736_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0737_
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1688980957
transform 1 0 16928 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0739_
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0740_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0741_
timestamp 1688980957
transform 1 0 17388 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0742_
timestamp 1688980957
transform 1 0 17296 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0743_
timestamp 1688980957
transform 1 0 17020 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1688980957
transform 1 0 17848 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0745_
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0746_
timestamp 1688980957
transform 1 0 17204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1688980957
transform 1 0 16836 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0748_
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0749_
timestamp 1688980957
transform 1 0 16744 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0750_
timestamp 1688980957
transform 1 0 17296 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0753_
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0754_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0755_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1688980957
transform 1 0 16560 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0757_
timestamp 1688980957
transform 1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1688980957
transform 1 0 15548 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0759_
timestamp 1688980957
transform 1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0760_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0761_
timestamp 1688980957
transform 1 0 14628 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0762_
timestamp 1688980957
transform 1 0 15824 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _0763_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0765_
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0767_
timestamp 1688980957
transform 1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0768_
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0769_
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0770_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0771_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0772_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0773_
timestamp 1688980957
transform 1 0 15824 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0774_
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0775_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0776_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0777_
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1688980957
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1688980957
transform 1 0 16560 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0781_
timestamp 1688980957
transform 1 0 13248 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0782_
timestamp 1688980957
transform 1 0 12512 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0784_
timestamp 1688980957
transform 1 0 15364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0785_
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0786_
timestamp 1688980957
transform 1 0 14720 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0787_
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0788_
timestamp 1688980957
transform 1 0 14812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0789_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0790_
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0791_
timestamp 1688980957
transform 1 0 14996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0792_
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0793_
timestamp 1688980957
transform 1 0 14720 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0794_
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_2  _0795_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1688980957
transform 1 0 12144 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0797_
timestamp 1688980957
transform 1 0 11592 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1688980957
transform 1 0 12696 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0799_
timestamp 1688980957
transform 1 0 11316 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0800_
timestamp 1688980957
transform 1 0 13524 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0802_
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0803_
timestamp 1688980957
transform 1 0 14168 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0804_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0805_
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _0806_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12144 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0807_
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0808_
timestamp 1688980957
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0809_
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0810_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0811_
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0812_
timestamp 1688980957
transform 1 0 20424 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0814_
timestamp 1688980957
transform 1 0 17848 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 1688980957
transform 1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0816_
timestamp 1688980957
transform 1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0817_
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0820_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0821_
timestamp 1688980957
transform 1 0 6992 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0822_
timestamp 1688980957
transform 1 0 8004 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0824_
timestamp 1688980957
transform 1 0 8372 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1688980957
transform 1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0826_
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1688980957
transform 1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0828_
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0829_
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0830_
timestamp 1688980957
transform 1 0 7176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 1688980957
transform 1 0 7268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0833_
timestamp 1688980957
transform 1 0 6440 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0835_
timestamp 1688980957
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0836_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0837_
timestamp 1688980957
transform 1 0 6072 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 1688980957
transform 1 0 7084 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 1688980957
transform 1 0 7912 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 1688980957
transform 1 0 8372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0841_
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 1688980957
transform 1 0 8188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0844_
timestamp 1688980957
transform 1 0 9384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0845_
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1688980957
transform 1 0 15732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0847_
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1688980957
transform 1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0849_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1688980957
transform 1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1688980957
transform 1 0 15824 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0852_
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0853_
timestamp 1688980957
transform 1 0 15088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0854_
timestamp 1688980957
transform 1 0 16192 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0858_
timestamp 1688980957
transform 1 0 12144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0860_
timestamp 1688980957
transform 1 0 16468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0861_
timestamp 1688980957
transform 1 0 17572 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0863_
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0864_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0865_
timestamp 1688980957
transform 1 0 15824 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0866_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16560 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0867_
timestamp 1688980957
transform 1 0 15916 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0868_
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0869_
timestamp 1688980957
transform 1 0 14168 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0870_
timestamp 1688980957
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0871_
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0872_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _0873_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _0874_
timestamp 1688980957
transform 1 0 15456 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0875_
timestamp 1688980957
transform 1 0 15088 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1688980957
transform 1 0 15272 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1688980957
transform 1 0 14904 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0879_
timestamp 1688980957
transform 1 0 15456 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0880_
timestamp 1688980957
transform 1 0 14904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0881_
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0883_
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0884_
timestamp 1688980957
transform 1 0 14260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0885_
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0886_
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0887_
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0888_
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0889_
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0890_
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0892_
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0893_
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0894_
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0895_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0896_
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0897_
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0898_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0899_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0900_
timestamp 1688980957
transform 1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0901_
timestamp 1688980957
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0902_
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0904_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0905_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0906_
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0907_
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0908_
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0910_
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0911_
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0912_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0913_
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0916_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0919_
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0920_
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0923_
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0925_
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0926_
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0927_
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0929_
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0930_
timestamp 1688980957
transform 1 0 15364 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0931_
timestamp 1688980957
transform 1 0 17388 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 1688980957
transform 1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0933_
timestamp 1688980957
transform 1 0 16744 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1688980957
transform 1 0 16836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0936_
timestamp 1688980957
transform 1 0 16192 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0937_
timestamp 1688980957
transform 1 0 17940 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0939_
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1688980957
transform 1 0 16008 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0941_
timestamp 1688980957
transform 1 0 15272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1688980957
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0943_
timestamp 1688980957
transform 1 0 16468 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0945_
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0946_
timestamp 1688980957
transform 1 0 15732 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0947_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0948_
timestamp 1688980957
transform 1 0 12788 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0949_
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0950_
timestamp 1688980957
transform 1 0 12696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0952_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0953_
timestamp 1688980957
transform 1 0 11684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1688980957
transform 1 0 20608 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 1688980957
transform 1 0 20884 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0960_
timestamp 1688980957
transform 1 0 18584 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0963_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1688980957
transform 1 0 21252 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0967_
timestamp 1688980957
transform 1 0 20700 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1688980957
transform 1 0 20240 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1688980957
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1688980957
transform 1 0 20148 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1688980957
transform 1 0 19872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp 1688980957
transform 1 0 20056 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1688980957
transform 1 0 20148 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0981_
timestamp 1688980957
transform 1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1688980957
transform 1 0 6164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1688980957
transform 1 0 7268 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp 1688980957
transform 1 0 9752 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1688980957
transform 1 0 20884 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1688980957
transform 1 0 21160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1688980957
transform 1 0 23460 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1688980957
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1688980957
transform 1 0 23368 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1688980957
transform 1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1688980957
transform 1 0 21896 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1688980957
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1688980957
transform 1 0 24380 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1688980957
transform 1 0 24472 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1688980957
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp 1688980957
transform 1 0 17020 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1688980957
transform 1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1020_
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1021_
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1022_
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1023_
timestamp 1688980957
transform 1 0 11776 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1024_
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1025_
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1026_
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1028_
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1031_
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1032_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1033_
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1034_
timestamp 1688980957
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1688980957
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1036_
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1688980957
transform 1 0 5704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1038_
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1040_
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1688980957
transform 1 0 6348 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1042_
timestamp 1688980957
transform 1 0 3128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1044_
timestamp 1688980957
transform 1 0 2576 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1046_
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1048_
timestamp 1688980957
transform 1 0 10488 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1050_
timestamp 1688980957
transform 1 0 4140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1052_
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1054_
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1056_
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1057_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1058_
timestamp 1688980957
transform 1 0 2944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1688980957
transform 1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1060_
timestamp 1688980957
transform 1 0 2760 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1688980957
transform 1 0 3312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1062_
timestamp 1688980957
transform 1 0 2208 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1063_
timestamp 1688980957
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1064_
timestamp 1688980957
transform 1 0 2392 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1688980957
transform 1 0 5152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1066_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1067_
timestamp 1688980957
transform 1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1068_
timestamp 1688980957
transform 1 0 20516 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1069_
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1070_
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1071_
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1072_
timestamp 1688980957
transform 1 0 21068 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1073_
timestamp 1688980957
transform 1 0 21620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1074_
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1688980957
transform 1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1076_
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1078_
timestamp 1688980957
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1079_
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1080_
timestamp 1688980957
transform 1 0 9936 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1082_
timestamp 1688980957
transform 1 0 9936 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 1688980957
transform 1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1084_
timestamp 1688980957
transform 1 0 4968 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1085_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1086_
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1087_
timestamp 1688980957
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1088_
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1688980957
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1090_
timestamp 1688980957
transform 1 0 6900 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1091_
timestamp 1688980957
transform 1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1092_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1093_
timestamp 1688980957
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1094_
timestamp 1688980957
transform 1 0 7544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1095_
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1096_
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1098_
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1099_
timestamp 1688980957
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1100_
timestamp 1688980957
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1688980957
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1102_
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1688980957
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1104_
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1106_
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1688980957
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1108_
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1688980957
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1110_
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1112_
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1113_
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1114_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1116_
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1117_
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1688980957
transform 1 0 17664 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1119_
timestamp 1688980957
transform 1 0 18216 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1120_
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1121_
timestamp 1688980957
transform 1 0 9384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1122_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1688980957
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1124_
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1126_
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1127_
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1128_
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1130_
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1131_
timestamp 1688980957
transform 1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1132_
timestamp 1688980957
transform 1 0 11776 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1134_
timestamp 1688980957
transform 1 0 12696 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1135_
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1136_
timestamp 1688980957
transform 1 0 12696 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1137_
timestamp 1688980957
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1138_
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1139_
timestamp 1688980957
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1140_
timestamp 1688980957
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1688980957
transform 1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1142_
timestamp 1688980957
transform 1 0 12696 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1144_
timestamp 1688980957
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1145_
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1146_
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1148_
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1688980957
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1150_
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1688980957
transform 1 0 14720 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1152_
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1688980957
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1154_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1156_
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1158_
timestamp 1688980957
transform 1 0 3864 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1160_
timestamp 1688980957
transform 1 0 4784 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1162_
timestamp 1688980957
transform 1 0 7912 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1688980957
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1164_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1165_
timestamp 1688980957
transform 1 0 10396 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1166_
timestamp 1688980957
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1167_
timestamp 1688980957
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1168_
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1170_
timestamp 1688980957
transform 1 0 14536 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1171_
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1172_
timestamp 1688980957
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1688980957
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1174_
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1688980957
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1178_
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1688980957
transform 1 0 18768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1180_
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1688980957
transform 1 0 18400 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1182_
timestamp 1688980957
transform 1 0 13156 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1184_
timestamp 1688980957
transform 1 0 12788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1185_
timestamp 1688980957
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1186_
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1187_
timestamp 1688980957
transform 1 0 13432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1688980957
transform 1 0 19320 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1189_
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1190_
timestamp 1688980957
transform 1 0 20976 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1688980957
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1192_
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1193_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1194_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1196_
timestamp 1688980957
transform 1 0 20148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1688980957
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1198_
timestamp 1688980957
transform 1 0 20332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1688980957
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1202_
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1204_
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1206_
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1208_
timestamp 1688980957
transform 1 0 20424 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1688980957
transform 1 0 20976 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1210_
timestamp 1688980957
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1211_
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1212_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1688980957
transform 1 0 19412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1214_
timestamp 1688980957
transform 1 0 19872 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1688980957
transform 1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1216_
timestamp 1688980957
transform 1 0 19688 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1688980957
transform 1 0 21160 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1218_
timestamp 1688980957
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1219_
timestamp 1688980957
transform 1 0 8280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1220_
timestamp 1688980957
transform 1 0 9200 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1221_
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1222_
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1688980957
transform 1 0 11776 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1224_
timestamp 1688980957
transform 1 0 19872 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1688980957
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1226_
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1228_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1229_
timestamp 1688980957
transform 1 0 18768 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1230_
timestamp 1688980957
transform 1 0 9844 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1688980957
transform 1 0 10396 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1232_
timestamp 1688980957
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1233_
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1234_
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1235_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1236_
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1688980957
transform 1 0 24932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1238_
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1688980957
transform 1 0 24472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1240_
timestamp 1688980957
transform 1 0 23368 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1241_
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1242_
timestamp 1688980957
transform 1 0 23552 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1243_
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1244_
timestamp 1688980957
transform 1 0 24932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1688980957
transform 1 0 24932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1246_
timestamp 1688980957
transform 1 0 23828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1247_
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1248_
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1688980957
transform 1 0 24656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1250_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1251_
timestamp 1688980957
transform 1 0 25300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1252_
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1254_
timestamp 1688980957
transform 1 0 17480 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1688980957
transform 1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1256_
timestamp 1688980957
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1258_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1259_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1688980957
transform 1 0 4324 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1688980957
transform 1 0 1656 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1688980957
transform 1 0 1564 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 1688980957
transform 1 0 11040 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1688980957
transform 1 0 3864 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1266_
timestamp 1688980957
transform 1 0 12420 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1267_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1688980957
transform 1 0 2668 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1269_
timestamp 1688980957
transform 1 0 2392 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1270_
timestamp 1688980957
transform 1 0 1840 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1271_
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 1688980957
transform 1 0 19596 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 1688980957
transform 1 0 20516 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1274_
timestamp 1688980957
transform 1 0 20884 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1275_
timestamp 1688980957
transform 1 0 20608 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1276_
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1277_
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1278_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1279_
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1280_
timestamp 1688980957
transform 1 0 5520 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 1688980957
transform 1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1282_
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1283_
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 1688980957
transform 1 0 6072 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 1688980957
transform 1 0 9016 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1688980957
transform 1 0 4232 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1291_
timestamp 1688980957
transform 1 0 14628 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1292_
timestamp 1688980957
transform 1 0 9108 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1293_
timestamp 1688980957
transform 1 0 8464 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1295_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1296_
timestamp 1688980957
transform 1 0 17204 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1297_
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1298_
timestamp 1688980957
transform 1 0 8372 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1299_
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1300_
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1301_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1303_
timestamp 1688980957
transform 1 0 13248 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1304_
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1305_
timestamp 1688980957
transform 1 0 11592 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1306_
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1307_
timestamp 1688980957
transform 1 0 13524 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1308_
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1309_
timestamp 1688980957
transform 1 0 14536 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1310_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1313_
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1314_
timestamp 1688980957
transform 1 0 3956 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1315_
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1316_
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1317_
timestamp 1688980957
transform 1 0 8740 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 1688980957
transform 1 0 10948 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1319_
timestamp 1688980957
transform 1 0 13892 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1320_
timestamp 1688980957
transform 1 0 16928 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1321_
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1322_
timestamp 1688980957
transform 1 0 15732 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1323_
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1324_
timestamp 1688980957
transform 1 0 17020 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1325_
timestamp 1688980957
transform 1 0 12420 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1328_
timestamp 1688980957
transform 1 0 20424 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 1688980957
transform 1 0 20884 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 1688980957
transform 1 0 20976 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1331_
timestamp 1688980957
transform 1 0 19872 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1332_
timestamp 1688980957
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1334_
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1335_
timestamp 1688980957
transform 1 0 19780 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 1688980957
transform 1 0 20516 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 1688980957
transform 1 0 19320 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 1688980957
transform 1 0 6440 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1342_
timestamp 1688980957
transform 1 0 8280 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 1688980957
transform 1 0 10764 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1344_
timestamp 1688980957
transform 1 0 20424 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1345_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 1688980957
transform 1 0 17848 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1347_
timestamp 1688980957
transform 1 0 8832 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1348_
timestamp 1688980957
transform 1 0 23460 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1349_
timestamp 1688980957
transform 1 0 23092 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1350_
timestamp 1688980957
transform 1 0 23736 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1351_
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1352_
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1688980957
transform 1 0 23092 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 1688980957
transform 1 0 23644 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1355_
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1356_
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 1688980957
transform 1 0 22632 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 1688980957
transform 1 0 16376 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1359_
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1688980957
transform 1 0 9568 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1688980957
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1688980957
transform 1 0 18216 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1688980957
transform 1 0 18216 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_12 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_44
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_51 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_90
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_104
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_164
timestamp 1688980957
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_178
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_231 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_244
timestamp 1688980957
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_24 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_36
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_101
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1688980957
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_136
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_160
timestamp 1688980957
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_178
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_190
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_202
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_214
timestamp 1688980957
transform 1 0 20792 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_234
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_246
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_12
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_24
timestamp 1688980957
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_33
timestamp 1688980957
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_106
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_182
timestamp 1688980957
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_244
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 1688980957
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_63
timestamp 1688980957
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_84
timestamp 1688980957
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_121
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_130
timestamp 1688980957
transform 1 0 13064 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_136
timestamp 1688980957
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_140
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 1688980957
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_175
timestamp 1688980957
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_185
timestamp 1688980957
transform 1 0 18124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_197
timestamp 1688980957
transform 1 0 19228 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_203
timestamp 1688980957
transform 1 0 19780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_231
timestamp 1688980957
transform 1 0 22356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_243
timestamp 1688980957
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_255
timestamp 1688980957
transform 1 0 24564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_263
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1688980957
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1688980957
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_119
timestamp 1688980957
transform 1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_123
timestamp 1688980957
transform 1 0 12420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_167
timestamp 1688980957
transform 1 0 16468 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_171
timestamp 1688980957
transform 1 0 16836 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_215
timestamp 1688980957
transform 1 0 20884 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_219
timestamp 1688980957
transform 1 0 21252 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_235
timestamp 1688980957
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 1688980957
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_261
timestamp 1688980957
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_30
timestamp 1688980957
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1688980957
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_133
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_143
timestamp 1688980957
transform 1 0 14260 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_185
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_206
timestamp 1688980957
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_231
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_243
timestamp 1688980957
transform 1 0 23460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_255
timestamp 1688980957
transform 1 0 24564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_62
timestamp 1688980957
transform 1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_113
timestamp 1688980957
transform 1 0 11500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_162
timestamp 1688980957
transform 1 0 16008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_184
timestamp 1688980957
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_188
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_203
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_235
timestamp 1688980957
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp 1688980957
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_82
timestamp 1688980957
transform 1 0 8648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_89
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_102
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_141
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_147
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_155
timestamp 1688980957
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_159
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_175
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_204
timestamp 1688980957
transform 1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_228
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_240
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_252
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_260
timestamp 1688980957
transform 1 0 25024 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_39
timestamp 1688980957
transform 1 0 4692 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_46
timestamp 1688980957
transform 1 0 5336 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_50
timestamp 1688980957
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_58
timestamp 1688980957
transform 1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 1688980957
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp 1688980957
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_173
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_179
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_19
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_41
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_49
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_140
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_190
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_195
timestamp 1688980957
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_207
timestamp 1688980957
transform 1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_215
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_234
timestamp 1688980957
transform 1 0 22632 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_246
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_258
timestamp 1688980957
transform 1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_24
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_39
timestamp 1688980957
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_51
timestamp 1688980957
transform 1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_92
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_104
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 1688980957
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_128
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_167
timestamp 1688980957
transform 1 0 16468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_184
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_213
timestamp 1688980957
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_234
timestamp 1688980957
transform 1 0 22632 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_259
timestamp 1688980957
transform 1 0 24932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_16
timestamp 1688980957
transform 1 0 2576 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_65
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_98
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_121
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_144
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_150
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_196
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1688980957
transform 1 0 19688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_215
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_228
timestamp 1688980957
transform 1 0 22080 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_240
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_19
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_38
timestamp 1688980957
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_99
timestamp 1688980957
transform 1 0 10212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_161
timestamp 1688980957
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_181
timestamp 1688980957
transform 1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_187
timestamp 1688980957
transform 1 0 18308 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_222
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_234
timestamp 1688980957
transform 1 0 22632 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_240
timestamp 1688980957
transform 1 0 23184 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_262
timestamp 1688980957
transform 1 0 25208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_30
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_76
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_104
timestamp 1688980957
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_108
timestamp 1688980957
transform 1 0 11040 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_144
timestamp 1688980957
transform 1 0 14352 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_184
timestamp 1688980957
transform 1 0 18032 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_206
timestamp 1688980957
transform 1 0 20056 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_218
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_233
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_51
timestamp 1688980957
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_63
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_67
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_92
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_104
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_110
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_172
timestamp 1688980957
transform 1 0 16928 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_206
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_224
timestamp 1688980957
transform 1 0 21712 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 1688980957
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_259
timestamp 1688980957
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_30
timestamp 1688980957
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_67
timestamp 1688980957
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_135
timestamp 1688980957
transform 1 0 13524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1688980957
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_195
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_228
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_234
timestamp 1688980957
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_17
timestamp 1688980957
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_69
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_73
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1688980957
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_111
timestamp 1688980957
transform 1 0 11316 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_123
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1688980957
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_168
timestamp 1688980957
transform 1 0 16560 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_205
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_220
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_232
timestamp 1688980957
transform 1 0 22448 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_239
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_259
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_6
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_62
timestamp 1688980957
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_66
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_70
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_74
timestamp 1688980957
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_89
timestamp 1688980957
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_122
timestamp 1688980957
transform 1 0 12328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_134
timestamp 1688980957
transform 1 0 13432 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_146
timestamp 1688980957
transform 1 0 14536 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_154
timestamp 1688980957
transform 1 0 15272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 1688980957
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_175
timestamp 1688980957
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_180
timestamp 1688980957
transform 1 0 17664 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_192
timestamp 1688980957
transform 1 0 18768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_204
timestamp 1688980957
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_212
timestamp 1688980957
transform 1 0 20608 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_234
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_246
timestamp 1688980957
transform 1 0 23736 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_252
timestamp 1688980957
transform 1 0 24288 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_262
timestamp 1688980957
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 1688980957
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_59
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_73
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1688980957
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_91
timestamp 1688980957
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_105
timestamp 1688980957
transform 1 0 10764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_151
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_163
timestamp 1688980957
transform 1 0 16100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_171
timestamp 1688980957
transform 1 0 16836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_202
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_231
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_239
timestamp 1688980957
transform 1 0 23092 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_38
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_42
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_82
timestamp 1688980957
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_94
timestamp 1688980957
transform 1 0 9752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_100
timestamp 1688980957
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_107
timestamp 1688980957
transform 1 0 10948 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1688980957
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1688980957
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_233
timestamp 1688980957
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_21
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_25
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_59
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_69
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_79
timestamp 1688980957
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_99
timestamp 1688980957
transform 1 0 10212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_107
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_118
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_162
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1688980957
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_200
timestamp 1688980957
transform 1 0 19504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_219
timestamp 1688980957
transform 1 0 21252 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_223
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_235
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_243
timestamp 1688980957
transform 1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_257
timestamp 1688980957
transform 1 0 24748 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 1688980957
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_18
timestamp 1688980957
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_31
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_50
timestamp 1688980957
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1688980957
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_160
timestamp 1688980957
transform 1 0 15824 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1688980957
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_6
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_24
timestamp 1688980957
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_74
timestamp 1688980957
transform 1 0 7912 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_96
timestamp 1688980957
transform 1 0 9936 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_102
timestamp 1688980957
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_124
timestamp 1688980957
transform 1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_175
timestamp 1688980957
transform 1 0 17204 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_183
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_192
timestamp 1688980957
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_231
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_235
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_243
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_257
timestamp 1688980957
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_30
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_60
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_71
timestamp 1688980957
transform 1 0 7636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_83
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_116
timestamp 1688980957
transform 1 0 11776 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_128
timestamp 1688980957
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_156
timestamp 1688980957
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_177
timestamp 1688980957
transform 1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 1688980957
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_215
timestamp 1688980957
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_235
timestamp 1688980957
transform 1 0 22724 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_265
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_24
timestamp 1688980957
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_93
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_99
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_104
timestamp 1688980957
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_127
timestamp 1688980957
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_131
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_155
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_217
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_13
timestamp 1688980957
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_36
timestamp 1688980957
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_48
timestamp 1688980957
transform 1 0 5520 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_73
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_95
timestamp 1688980957
transform 1 0 9844 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_122
timestamp 1688980957
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_143
timestamp 1688980957
transform 1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_151
timestamp 1688980957
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_210
timestamp 1688980957
transform 1 0 20424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1688980957
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_231
timestamp 1688980957
transform 1 0 22356 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_235
timestamp 1688980957
transform 1 0 22724 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_265
timestamp 1688980957
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_56
timestamp 1688980957
transform 1 0 6256 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_60
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_72
timestamp 1688980957
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_128
timestamp 1688980957
transform 1 0 12880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_159
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_171
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_179
timestamp 1688980957
transform 1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_190
timestamp 1688980957
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_241
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_264
timestamp 1688980957
transform 1 0 25392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_33
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_61
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_88
timestamp 1688980957
transform 1 0 9200 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_100
timestamp 1688980957
transform 1 0 10304 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_134
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_162
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_173
timestamp 1688980957
transform 1 0 17020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_185
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_197
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_204
timestamp 1688980957
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 1688980957
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_234
timestamp 1688980957
transform 1 0 22632 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_245
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_259
timestamp 1688980957
transform 1 0 24932 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1688980957
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_35
timestamp 1688980957
transform 1 0 4324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_43
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_106
timestamp 1688980957
transform 1 0 10856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_114
timestamp 1688980957
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_206
timestamp 1688980957
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_210
timestamp 1688980957
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_262
timestamp 1688980957
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_9
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_14
timestamp 1688980957
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_26
timestamp 1688980957
transform 1 0 3496 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_34
timestamp 1688980957
transform 1 0 4232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_63
timestamp 1688980957
transform 1 0 6900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_68
timestamp 1688980957
transform 1 0 7360 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_86
timestamp 1688980957
transform 1 0 9016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_99
timestamp 1688980957
transform 1 0 10212 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_103
timestamp 1688980957
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_134
timestamp 1688980957
transform 1 0 13432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_178
timestamp 1688980957
transform 1 0 17480 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_185
timestamp 1688980957
transform 1 0 18124 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_206
timestamp 1688980957
transform 1 0 20056 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_218
timestamp 1688980957
transform 1 0 21160 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_234
timestamp 1688980957
transform 1 0 22632 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_238
timestamp 1688980957
transform 1 0 23000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_260
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_38
timestamp 1688980957
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_50
timestamp 1688980957
transform 1 0 5704 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_59
timestamp 1688980957
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_71
timestamp 1688980957
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_119
timestamp 1688980957
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_131
timestamp 1688980957
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_183
timestamp 1688980957
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_203
timestamp 1688980957
transform 1 0 19780 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_211
timestamp 1688980957
transform 1 0 20516 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_12
timestamp 1688980957
transform 1 0 2208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_37
timestamp 1688980957
transform 1 0 4508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1688980957
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_92
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_100
timestamp 1688980957
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_172
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_180
timestamp 1688980957
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_232
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_263
timestamp 1688980957
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_47
timestamp 1688980957
transform 1 0 5428 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_74
timestamp 1688980957
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_173
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_181
timestamp 1688980957
transform 1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_187
timestamp 1688980957
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_206
timestamp 1688980957
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_210
timestamp 1688980957
transform 1 0 20424 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_238
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_242
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_256
timestamp 1688980957
transform 1 0 24656 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_32
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_44
timestamp 1688980957
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_74
timestamp 1688980957
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_78
timestamp 1688980957
transform 1 0 8280 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_103
timestamp 1688980957
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_130
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_142
timestamp 1688980957
transform 1 0 14168 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_154
timestamp 1688980957
transform 1 0 15272 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_187
timestamp 1688980957
transform 1 0 18308 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_192
timestamp 1688980957
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_208
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_213
timestamp 1688980957
transform 1 0 20700 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_219
timestamp 1688980957
transform 1 0 21252 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_234
timestamp 1688980957
transform 1 0 22632 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_242
timestamp 1688980957
transform 1 0 23368 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_247
timestamp 1688980957
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_259
timestamp 1688980957
transform 1 0 24932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_265
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_6
timestamp 1688980957
transform 1 0 1656 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_50
timestamp 1688980957
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_62
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_74
timestamp 1688980957
transform 1 0 7912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_80
timestamp 1688980957
transform 1 0 8464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_105
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_116
timestamp 1688980957
transform 1 0 11776 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_123
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_150
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_178
timestamp 1688980957
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_190
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_235
timestamp 1688980957
transform 1 0 22724 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1688980957
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_261
timestamp 1688980957
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_9
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_34
timestamp 1688980957
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_70
timestamp 1688980957
transform 1 0 7544 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_103
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_131
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_156
timestamp 1688980957
transform 1 0 15456 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_164
timestamp 1688980957
transform 1 0 16192 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_183
timestamp 1688980957
transform 1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_189
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_215
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_252
timestamp 1688980957
transform 1 0 24288 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_264
timestamp 1688980957
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_7
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_46
timestamp 1688980957
transform 1 0 5336 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_56
timestamp 1688980957
transform 1 0 6256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_68
timestamp 1688980957
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_112
timestamp 1688980957
transform 1 0 11408 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_125
timestamp 1688980957
transform 1 0 12604 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_186
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_220
timestamp 1688980957
transform 1 0 21344 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_232
timestamp 1688980957
transform 1 0 22448 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_244
timestamp 1688980957
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_261
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_9
timestamp 1688980957
transform 1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_13
timestamp 1688980957
transform 1 0 2300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_17
timestamp 1688980957
transform 1 0 2668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_82
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_100
timestamp 1688980957
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_146
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_152
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_160
timestamp 1688980957
transform 1 0 15824 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_187
timestamp 1688980957
transform 1 0 18308 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_68
timestamp 1688980957
transform 1 0 7360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_80
timestamp 1688980957
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_108
timestamp 1688980957
transform 1 0 11040 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_128
timestamp 1688980957
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_144
timestamp 1688980957
transform 1 0 14352 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_164
timestamp 1688980957
transform 1 0 16192 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_181
timestamp 1688980957
transform 1 0 17756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_203
timestamp 1688980957
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_210
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_6
timestamp 1688980957
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_18
timestamp 1688980957
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_30
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_42
timestamp 1688980957
transform 1 0 4968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_52
timestamp 1688980957
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_64
timestamp 1688980957
transform 1 0 6992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_76
timestamp 1688980957
transform 1 0 8096 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_80
timestamp 1688980957
transform 1 0 8464 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_88
timestamp 1688980957
transform 1 0 9200 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_101
timestamp 1688980957
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_122
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_134
timestamp 1688980957
transform 1 0 13432 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_140
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_152
timestamp 1688980957
transform 1 0 15088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_158
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_174
timestamp 1688980957
transform 1 0 17112 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_186
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_198
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_206
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_210
timestamp 1688980957
transform 1 0 20424 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_214
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_245
timestamp 1688980957
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_257
timestamp 1688980957
transform 1 0 24748 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_7
timestamp 1688980957
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_19
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_73
timestamp 1688980957
transform 1 0 7820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_79
timestamp 1688980957
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_110
timestamp 1688980957
transform 1 0 11224 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_131
timestamp 1688980957
transform 1 0 13156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_152
timestamp 1688980957
transform 1 0 15088 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_156
timestamp 1688980957
transform 1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_180
timestamp 1688980957
transform 1 0 17664 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_192
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_201
timestamp 1688980957
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_208
timestamp 1688980957
transform 1 0 20240 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_215
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_224
timestamp 1688980957
transform 1 0 21712 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_236
timestamp 1688980957
transform 1 0 22816 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_261
timestamp 1688980957
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_66
timestamp 1688980957
transform 1 0 7176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_124
timestamp 1688980957
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_187
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_195
timestamp 1688980957
transform 1 0 19044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_265
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_12
timestamp 1688980957
transform 1 0 2208 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_24
timestamp 1688980957
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_103
timestamp 1688980957
transform 1 0 10580 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_125
timestamp 1688980957
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_132
timestamp 1688980957
transform 1 0 13248 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_136
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_191
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_203
timestamp 1688980957
transform 1 0 19780 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_230
timestamp 1688980957
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_242
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_248
timestamp 1688980957
transform 1 0 23920 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_25
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_37
timestamp 1688980957
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_49
timestamp 1688980957
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_131
timestamp 1688980957
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_143
timestamp 1688980957
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_155
timestamp 1688980957
transform 1 0 15364 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_163
timestamp 1688980957
transform 1 0 16100 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_177
timestamp 1688980957
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_202
timestamp 1688980957
transform 1 0 19688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_210
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_245
timestamp 1688980957
transform 1 0 23644 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_9
timestamp 1688980957
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_16
timestamp 1688980957
transform 1 0 2576 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_32
timestamp 1688980957
transform 1 0 4048 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_44
timestamp 1688980957
transform 1 0 5152 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_48
timestamp 1688980957
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_55
timestamp 1688980957
transform 1 0 6164 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_57
timestamp 1688980957
transform 1 0 6348 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_62
timestamp 1688980957
transform 1 0 6808 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_72
timestamp 1688980957
transform 1 0 7728 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_105
timestamp 1688980957
transform 1 0 10764 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_113
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_132
timestamp 1688980957
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_156
timestamp 1688980957
transform 1 0 15456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_160
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_169
timestamp 1688980957
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_181
timestamp 1688980957
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_188
timestamp 1688980957
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_203
timestamp 1688980957
transform 1 0 19780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_219
timestamp 1688980957
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_223
timestamp 1688980957
transform 1 0 21620 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_234
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_244
timestamp 1688980957
transform 1 0 23552 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 10120 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 12696 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 8096 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 16100 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 19688 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 3772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 21712 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 21988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 15548 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 24748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 25300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 25300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 22356 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 25300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 9476 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 25300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 25024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 12328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 12972 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 9752 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 18124 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 25024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1688980957
transform 1 0 2668 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1688980957
transform 1 0 24564 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 23736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 25300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1688980957
transform 1 0 24656 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 24932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  max_cap133
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 14260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 21804 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 2024 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 10856 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1688980957
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 25024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 24104 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1688980957
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1688980957
transform 1 0 25208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 25024 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform 1 0 25208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 25024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 11684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 24656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 25208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 24472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform 1 0 24656 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 7176 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 20700 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 14904 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 1748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1688980957
transform 1 0 25208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 15640 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 20056 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 2300 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 6256 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 16560 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 21712 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
<< labels >>
flabel metal3 s 26237 23128 27037 23248 0 FreeSans 480 0 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 15474 28381 15530 29181 0 FreeSans 224 90 0 0 A[10]
port 1 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 A[11]
port 2 nsew signal input
flabel metal3 s 26237 688 27037 808 0 FreeSans 480 0 0 0 A[12]
port 3 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 A[13]
port 4 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 A[14]
port 5 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 A[15]
port 6 nsew signal input
flabel metal3 s 26237 26528 27037 26648 0 FreeSans 480 0 0 0 A[16]
port 7 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 A[17]
port 8 nsew signal input
flabel metal2 s 17406 28381 17462 29181 0 FreeSans 224 90 0 0 A[18]
port 9 nsew signal input
flabel metal2 s 3238 28381 3294 29181 0 FreeSans 224 90 0 0 A[19]
port 10 nsew signal input
flabel metal3 s 26237 8168 27037 8288 0 FreeSans 480 0 0 0 A[1]
port 11 nsew signal input
flabel metal3 s 26237 21768 27037 21888 0 FreeSans 480 0 0 0 A[20]
port 12 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 A[21]
port 13 nsew signal input
flabel metal2 s 25778 28381 25834 29181 0 FreeSans 224 90 0 0 A[22]
port 14 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 A[23]
port 15 nsew signal input
flabel metal3 s 26237 22448 27037 22568 0 FreeSans 480 0 0 0 A[24]
port 16 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 A[25]
port 17 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 A[26]
port 18 nsew signal input
flabel metal3 s 26237 10888 27037 11008 0 FreeSans 480 0 0 0 A[27]
port 19 nsew signal input
flabel metal3 s 26237 8 27037 128 0 FreeSans 480 0 0 0 A[28]
port 20 nsew signal input
flabel metal3 s 26237 3408 27037 3528 0 FreeSans 480 0 0 0 A[29]
port 21 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 A[2]
port 22 nsew signal input
flabel metal2 s 5814 28381 5870 29181 0 FreeSans 224 90 0 0 A[30]
port 23 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 A[31]
port 24 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 A[3]
port 25 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 A[4]
port 26 nsew signal input
flabel metal2 s 21914 28381 21970 29181 0 FreeSans 224 90 0 0 A[5]
port 27 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 A[6]
port 28 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 A[7]
port 29 nsew signal input
flabel metal3 s 26237 18368 27037 18488 0 FreeSans 480 0 0 0 A[8]
port 30 nsew signal input
flabel metal2 s 9034 28381 9090 29181 0 FreeSans 224 90 0 0 A[9]
port 31 nsew signal input
flabel metal2 s 5170 28381 5226 29181 0 FreeSans 224 90 0 0 B[0]
port 32 nsew signal input
flabel metal2 s 23202 28381 23258 29181 0 FreeSans 224 90 0 0 B[10]
port 33 nsew signal input
flabel metal3 s 26237 16328 27037 16448 0 FreeSans 480 0 0 0 B[11]
port 34 nsew signal input
flabel metal3 s 26237 17008 27037 17128 0 FreeSans 480 0 0 0 B[12]
port 35 nsew signal input
flabel metal2 s 12254 28381 12310 29181 0 FreeSans 224 90 0 0 B[13]
port 36 nsew signal input
flabel metal2 s 12898 28381 12954 29181 0 FreeSans 224 90 0 0 B[14]
port 37 nsew signal input
flabel metal2 s 9678 28381 9734 29181 0 FreeSans 224 90 0 0 B[15]
port 38 nsew signal input
flabel metal2 s 18050 28381 18106 29181 0 FreeSans 224 90 0 0 B[16]
port 39 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 B[17]
port 40 nsew signal input
flabel metal2 s 662 28381 718 29181 0 FreeSans 224 90 0 0 B[18]
port 41 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 B[19]
port 42 nsew signal input
flabel metal3 s 26237 12248 27037 12368 0 FreeSans 480 0 0 0 B[1]
port 43 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 B[20]
port 44 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 B[21]
port 45 nsew signal input
flabel metal3 s 26237 7488 27037 7608 0 FreeSans 480 0 0 0 B[22]
port 46 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 B[23]
port 47 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 B[24]
port 48 nsew signal input
flabel metal2 s 2594 28381 2650 29181 0 FreeSans 224 90 0 0 B[25]
port 49 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 B[26]
port 50 nsew signal input
flabel metal2 s 24490 28381 24546 29181 0 FreeSans 224 90 0 0 B[27]
port 51 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 B[28]
port 52 nsew signal input
flabel metal3 s 26237 28568 27037 28688 0 FreeSans 480 0 0 0 B[29]
port 53 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 B[2]
port 54 nsew signal input
flabel metal3 s 26237 20408 27037 20528 0 FreeSans 480 0 0 0 B[30]
port 55 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 B[31]
port 56 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 B[3]
port 57 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 B[4]
port 58 nsew signal input
flabel metal2 s 26422 28381 26478 29181 0 FreeSans 224 90 0 0 B[5]
port 59 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 B[6]
port 60 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 B[7]
port 61 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 B[8]
port 62 nsew signal input
flabel metal2 s 6458 28381 6514 29181 0 FreeSans 224 90 0 0 B[9]
port 63 nsew signal input
flabel metal2 s 14186 28381 14242 29181 0 FreeSans 224 90 0 0 D[0]
port 64 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 D[10]
port 65 nsew signal tristate
flabel metal2 s 21270 28381 21326 29181 0 FreeSans 224 90 0 0 D[11]
port 66 nsew signal tristate
flabel metal2 s 1950 28381 2006 29181 0 FreeSans 224 90 0 0 D[12]
port 67 nsew signal tristate
flabel metal2 s 8390 28381 8446 29181 0 FreeSans 224 90 0 0 D[13]
port 68 nsew signal tristate
flabel metal2 s 10966 28381 11022 29181 0 FreeSans 224 90 0 0 D[14]
port 69 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 D[15]
port 70 nsew signal tristate
flabel metal3 s 26237 12928 27037 13048 0 FreeSans 480 0 0 0 D[16]
port 71 nsew signal tristate
flabel metal3 s 26237 9528 27037 9648 0 FreeSans 480 0 0 0 D[17]
port 72 nsew signal tristate
flabel metal3 s 26237 25848 27037 25968 0 FreeSans 480 0 0 0 D[18]
port 73 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 D[19]
port 74 nsew signal tristate
flabel metal3 s 26237 1368 27037 1488 0 FreeSans 480 0 0 0 D[1]
port 75 nsew signal tristate
flabel metal3 s 26237 10208 27037 10328 0 FreeSans 480 0 0 0 D[20]
port 76 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 D[21]
port 77 nsew signal tristate
flabel metal3 s 26237 6128 27037 6248 0 FreeSans 480 0 0 0 D[22]
port 78 nsew signal tristate
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 D[23]
port 79 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 D[24]
port 80 nsew signal tristate
flabel metal3 s 26237 14288 27037 14408 0 FreeSans 480 0 0 0 D[25]
port 81 nsew signal tristate
flabel metal3 s 26237 27888 27037 28008 0 FreeSans 480 0 0 0 D[26]
port 82 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 D[27]
port 83 nsew signal tristate
flabel metal3 s 26237 4088 27037 4208 0 FreeSans 480 0 0 0 D[28]
port 84 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 D[29]
port 85 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 D[2]
port 86 nsew signal tristate
flabel metal2 s 11610 28381 11666 29181 0 FreeSans 224 90 0 0 D[30]
port 87 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 D[31]
port 88 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 D[3]
port 89 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 D[4]
port 90 nsew signal tristate
flabel metal3 s 26237 2728 27037 2848 0 FreeSans 480 0 0 0 D[5]
port 91 nsew signal tristate
flabel metal3 s 26237 19728 27037 19848 0 FreeSans 480 0 0 0 D[6]
port 92 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 D[7]
port 93 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 D[8]
port 94 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 D[9]
port 95 nsew signal tristate
flabel metal3 s 26237 6808 27037 6928 0 FreeSans 480 0 0 0 R[0]
port 96 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 R[10]
port 97 nsew signal tristate
flabel metal3 s 26237 15648 27037 15768 0 FreeSans 480 0 0 0 R[11]
port 98 nsew signal tristate
flabel metal3 s 26237 23808 27037 23928 0 FreeSans 480 0 0 0 R[12]
port 99 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 R[13]
port 100 nsew signal tristate
flabel metal3 s 26237 25168 27037 25288 0 FreeSans 480 0 0 0 R[14]
port 101 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 R[15]
port 102 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 R[16]
port 103 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 R[17]
port 104 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 R[18]
port 105 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 R[19]
port 106 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 R[1]
port 107 nsew signal tristate
flabel metal2 s 7102 28381 7158 29181 0 FreeSans 224 90 0 0 R[20]
port 108 nsew signal tristate
flabel metal2 s 16762 28381 16818 29181 0 FreeSans 224 90 0 0 R[21]
port 109 nsew signal tristate
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 R[22]
port 110 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 R[23]
port 111 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 R[24]
port 112 nsew signal tristate
flabel metal2 s 20626 28381 20682 29181 0 FreeSans 224 90 0 0 R[25]
port 113 nsew signal tristate
flabel metal2 s 14830 28381 14886 29181 0 FreeSans 224 90 0 0 R[26]
port 114 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 R[27]
port 115 nsew signal tristate
flabel metal2 s 23846 28381 23902 29181 0 FreeSans 224 90 0 0 R[28]
port 116 nsew signal tristate
flabel metal3 s 26237 4768 27037 4888 0 FreeSans 480 0 0 0 R[29]
port 117 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 R[2]
port 118 nsew signal tristate
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 R[30]
port 119 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 R[31]
port 120 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 R[3]
port 121 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 R[4]
port 122 nsew signal tristate
flabel metal3 s 26237 19048 27037 19168 0 FreeSans 480 0 0 0 R[5]
port 123 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 R[6]
port 124 nsew signal tristate
flabel metal2 s 19982 28381 20038 29181 0 FreeSans 224 90 0 0 R[7]
port 125 nsew signal tristate
flabel metal2 s 18694 28381 18750 29181 0 FreeSans 224 90 0 0 R[8]
port 126 nsew signal tristate
flabel metal2 s 18 28381 74 29181 0 FreeSans 224 90 0 0 R[9]
port 127 nsew signal tristate
flabel metal4 s 4697 2128 5017 26704 0 FreeSans 1920 90 0 0 VGND
port 128 nsew ground bidirectional
flabel metal4 s 10884 2128 11204 26704 0 FreeSans 1920 90 0 0 VGND
port 128 nsew ground bidirectional
flabel metal4 s 17071 2128 17391 26704 0 FreeSans 1920 90 0 0 VGND
port 128 nsew ground bidirectional
flabel metal4 s 23258 2128 23578 26704 0 FreeSans 1920 90 0 0 VGND
port 128 nsew ground bidirectional
flabel metal5 s 1056 5736 25900 6056 0 FreeSans 2560 0 0 0 VGND
port 128 nsew ground bidirectional
flabel metal5 s 1056 11856 25900 12176 0 FreeSans 2560 0 0 0 VGND
port 128 nsew ground bidirectional
flabel metal5 s 1056 17976 25900 18296 0 FreeSans 2560 0 0 0 VGND
port 128 nsew ground bidirectional
flabel metal5 s 1056 24096 25900 24416 0 FreeSans 2560 0 0 0 VGND
port 128 nsew ground bidirectional
flabel metal4 s 4037 2128 4357 26704 0 FreeSans 1920 90 0 0 VPWR
port 129 nsew power bidirectional
flabel metal4 s 10224 2128 10544 26704 0 FreeSans 1920 90 0 0 VPWR
port 129 nsew power bidirectional
flabel metal4 s 16411 2128 16731 26704 0 FreeSans 1920 90 0 0 VPWR
port 129 nsew power bidirectional
flabel metal4 s 22598 2128 22918 26704 0 FreeSans 1920 90 0 0 VPWR
port 129 nsew power bidirectional
flabel metal5 s 1056 5076 25900 5396 0 FreeSans 2560 0 0 0 VPWR
port 129 nsew power bidirectional
flabel metal5 s 1056 11196 25900 11516 0 FreeSans 2560 0 0 0 VPWR
port 129 nsew power bidirectional
flabel metal5 s 1056 17316 25900 17636 0 FreeSans 2560 0 0 0 VPWR
port 129 nsew power bidirectional
flabel metal5 s 1056 23436 25900 23756 0 FreeSans 2560 0 0 0 VPWR
port 129 nsew power bidirectional
flabel metal2 s 3882 28381 3938 29181 0 FreeSans 224 90 0 0 clk
port 130 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 err
port 131 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 ok
port 132 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 reset
port 133 nsew signal input
flabel metal3 s 26237 13608 27037 13728 0 FreeSans 480 0 0 0 start
port 134 nsew signal input
rlabel metal1 13478 26112 13478 26112 0 VGND
rlabel metal1 13478 26656 13478 26656 0 VPWR
rlabel metal1 25576 23698 25576 23698 0 A[0]
rlabel metal1 15640 26350 15640 26350 0 A[10]
rlabel metal2 23874 1027 23874 1027 0 A[11]
rlabel via2 25093 884 25093 884 0 A[12]
rlabel metal2 2806 7123 2806 7123 0 A[13]
rlabel metal3 820 4828 820 4828 0 A[14]
rlabel metal2 7774 1588 7774 1588 0 A[15]
rlabel metal1 23230 26316 23230 26316 0 A[16]
rlabel metal3 1050 23188 1050 23188 0 A[17]
rlabel metal1 17572 26350 17572 26350 0 A[18]
rlabel metal1 3634 26350 3634 26350 0 A[19]
rlabel metal1 25760 7854 25760 7854 0 A[1]
rlabel metal1 25530 21964 25530 21964 0 A[20]
rlabel metal3 866 25228 866 25228 0 A[21]
rlabel metal1 25024 25330 25024 25330 0 A[22]
rlabel metal2 12282 1588 12282 1588 0 A[23]
rlabel metal1 25530 22576 25530 22576 0 A[24]
rlabel metal2 7130 1588 7130 1588 0 A[25]
rlabel metal3 820 17068 820 17068 0 A[26]
rlabel metal1 25760 11118 25760 11118 0 A[27]
rlabel metal3 26136 68 26136 68 0 A[28]
rlabel metal1 25760 3502 25760 3502 0 A[29]
rlabel metal2 16790 1027 16790 1027 0 A[2]
rlabel metal1 5888 26350 5888 26350 0 A[30]
rlabel metal2 10994 1027 10994 1027 0 A[31]
rlabel metal2 25806 1146 25806 1146 0 A[3]
rlabel metal3 1050 20468 1050 20468 0 A[4]
rlabel metal1 22264 26350 22264 26350 0 A[5]
rlabel metal3 820 4148 820 4148 0 A[6]
rlabel metal3 820 11628 820 11628 0 A[7]
rlabel metal1 25530 18292 25530 18292 0 A[8]
rlabel metal1 9430 26350 9430 26350 0 A[9]
rlabel metal1 5244 26350 5244 26350 0 B[0]
rlabel metal1 23322 26384 23322 26384 0 B[10]
rlabel metal1 25760 17170 25760 17170 0 B[11]
rlabel metal1 25070 17136 25070 17136 0 B[12]
rlabel metal1 12328 26350 12328 26350 0 B[13]
rlabel metal1 12972 26350 12972 26350 0 B[14]
rlabel metal1 9752 26350 9752 26350 0 B[15]
rlabel metal1 18124 26350 18124 26350 0 B[16]
rlabel metal3 820 14348 820 14348 0 B[17]
rlabel metal2 690 27210 690 27210 0 B[18]
rlabel metal2 22586 959 22586 959 0 B[19]
rlabel metal1 25714 12818 25714 12818 0 B[1]
rlabel metal2 9062 1588 9062 1588 0 B[20]
rlabel metal2 13570 1588 13570 1588 0 B[21]
rlabel metal1 25070 7820 25070 7820 0 B[22]
rlabel metal2 6486 1588 6486 1588 0 B[23]
rlabel metal2 690 1860 690 1860 0 B[24]
rlabel metal2 2714 27455 2714 27455 0 B[25]
rlabel metal2 20010 1027 20010 1027 0 B[26]
rlabel metal2 24610 27455 24610 27455 0 B[27]
rlabel metal3 843 19108 843 19108 0 B[28]
rlabel metal1 23368 25874 23368 25874 0 B[29]
rlabel metal2 19366 1027 19366 1027 0 B[2]
rlabel metal1 25668 20910 25668 20910 0 B[30]
rlabel metal3 1050 13668 1050 13668 0 B[31]
rlabel metal2 10350 1588 10350 1588 0 B[3]
rlabel metal2 3910 1027 3910 1027 0 B[4]
rlabel metal1 24702 25772 24702 25772 0 B[5]
rlabel metal2 2898 26231 2898 26231 0 B[6]
rlabel metal3 866 3468 866 3468 0 B[7]
rlabel metal3 751 16388 751 16388 0 B[8]
rlabel metal1 6532 26350 6532 26350 0 B[9]
rlabel metal2 14490 27523 14490 27523 0 D[0]
rlabel metal3 751 19788 751 19788 0 D[10]
rlabel metal1 21666 26214 21666 26214 0 D[11]
rlabel metal2 2254 27523 2254 27523 0 D[12]
rlabel metal1 8786 26554 8786 26554 0 D[13]
rlabel metal2 11086 26979 11086 26979 0 D[14]
rlabel metal3 820 21148 820 21148 0 D[15]
rlabel metal2 25438 13073 25438 13073 0 D[16]
rlabel metal1 25714 9894 25714 9894 0 D[17]
rlabel metal1 24978 25874 24978 25874 0 D[18]
rlabel metal1 2346 2890 2346 2890 0 D[19]
rlabel metal3 25538 1428 25538 1428 0 D[1]
rlabel metal2 25438 10353 25438 10353 0 D[20]
rlabel metal3 1142 5508 1142 5508 0 D[21]
rlabel via2 25438 6171 25438 6171 0 D[22]
rlabel metal2 1610 27591 1610 27591 0 D[23]
rlabel metal3 820 15708 820 15708 0 D[24]
rlabel metal1 25714 14586 25714 14586 0 D[25]
rlabel metal1 25484 25466 25484 25466 0 D[26]
rlabel metal3 1142 10948 1142 10948 0 D[27]
rlabel metal2 25438 4301 25438 4301 0 D[28]
rlabel metal2 16146 823 16146 823 0 D[29]
rlabel metal2 25162 1520 25162 1520 0 D[2]
rlabel metal1 11776 26554 11776 26554 0 D[30]
rlabel metal2 21298 823 21298 823 0 D[31]
rlabel metal2 3266 959 3266 959 0 D[3]
rlabel metal3 820 10268 820 10268 0 D[4]
rlabel metal1 25116 2822 25116 2822 0 D[5]
rlabel metal1 25714 20026 25714 20026 0 D[6]
rlabel metal3 1740 748 1740 748 0 D[7]
rlabel metal2 21942 1690 21942 1690 0 D[8]
rlabel metal3 751 17748 751 17748 0 D[9]
rlabel metal1 25714 7174 25714 7174 0 R[0]
rlabel metal3 1004 1428 1004 1428 0 R[10]
rlabel via2 25438 15691 25438 15691 0 R[11]
rlabel metal2 25438 23953 25438 23953 0 R[12]
rlabel metal2 24518 823 24518 823 0 R[13]
rlabel metal2 24886 25347 24886 25347 0 R[14]
rlabel metal2 14858 959 14858 959 0 R[15]
rlabel metal3 820 12988 820 12988 0 R[16]
rlabel metal3 820 9588 820 9588 0 R[17]
rlabel metal1 828 2822 828 2822 0 R[18]
rlabel metal2 18078 1520 18078 1520 0 R[19]
rlabel metal1 1518 25466 1518 25466 0 R[1]
rlabel metal2 7406 27523 7406 27523 0 R[20]
rlabel metal1 16928 26554 16928 26554 0 R[21]
rlabel metal3 820 22508 820 22508 0 R[22]
rlabel metal2 4554 959 4554 959 0 R[23]
rlabel metal2 1334 959 1334 959 0 R[24]
rlabel metal1 20838 26554 20838 26554 0 R[25]
rlabel metal1 14996 26214 14996 26214 0 R[26]
rlabel metal2 12926 1520 12926 1520 0 R[27]
rlabel metal2 23966 27523 23966 27523 0 R[28]
rlabel metal2 25438 4913 25438 4913 0 R[29]
rlabel metal3 866 25908 866 25908 0 R[2]
rlabel metal3 1188 8228 1188 8228 0 R[30]
rlabel metal2 5198 959 5198 959 0 R[31]
rlabel metal2 9706 1520 9706 1520 0 R[3]
rlabel metal3 1142 2108 1142 2108 0 R[4]
rlabel metal2 25438 19023 25438 19023 0 R[5]
rlabel metal2 15502 1520 15502 1520 0 R[6]
rlabel metal1 20148 26554 20148 26554 0 R[7]
rlabel metal1 19274 26554 19274 26554 0 R[8]
rlabel metal1 1288 25670 1288 25670 0 R[9]
rlabel metal2 5750 15640 5750 15640 0 _0000_
rlabel metal2 6026 17000 6026 17000 0 _0001_
rlabel metal2 6394 17544 6394 17544 0 _0002_
rlabel metal2 2254 17442 2254 17442 0 _0003_
rlabel metal1 3135 16490 3135 16490 0 _0004_
rlabel metal1 3036 14586 3036 14586 0 _0005_
rlabel metal2 12466 16762 12466 16762 0 _0006_
rlabel metal1 5435 12206 5435 12206 0 _0007_
rlabel metal1 12604 15674 12604 15674 0 _0008_
rlabel metal2 11546 14552 11546 14552 0 _0009_
rlabel metal2 3542 19822 3542 19822 0 _0010_
rlabel metal2 3358 21352 3358 21352 0 _0011_
rlabel metal2 2162 21794 2162 21794 0 _0012_
rlabel metal1 4186 19958 4186 19958 0 _0013_
rlabel metal1 20095 19414 20095 19414 0 _0014_
rlabel metal2 21298 17816 21298 17816 0 _0015_
rlabel metal1 21567 20842 21567 20842 0 _0016_
rlabel metal2 21574 19176 21574 19176 0 _0017_
rlabel metal1 19458 18938 19458 18938 0 _0018_
rlabel metal2 12834 20162 12834 20162 0 _0019_
rlabel metal2 12466 17816 12466 17816 0 _0020_
rlabel metal2 10626 18258 10626 18258 0 _0021_
rlabel metal2 6394 14178 6394 14178 0 _0022_
rlabel metal1 4646 11832 4646 11832 0 _0023_
rlabel metal2 4646 13022 4646 13022 0 _0024_
rlabel metal1 7038 13498 7038 13498 0 _0025_
rlabel metal1 7176 3162 7176 3162 0 _0026_
rlabel metal1 10212 3366 10212 3366 0 _0027_
rlabel metal2 10350 4318 10350 4318 0 _0028_
rlabel metal1 5934 2890 5934 2890 0 _0029_
rlabel metal2 12466 5406 12466 5406 0 _0030_
rlabel metal2 12374 6562 12374 6562 0 _0031_
rlabel metal2 19366 6766 19366 6766 0 _0032_
rlabel metal2 15594 7650 15594 7650 0 _0033_
rlabel metal1 10817 11118 10817 11118 0 _0034_
rlabel metal1 10035 13974 10035 13974 0 _0035_
rlabel metal1 12144 11594 12144 11594 0 _0036_
rlabel metal2 19826 15266 19826 15266 0 _0037_
rlabel metal2 18262 15640 18262 15640 0 _0038_
rlabel metal1 9384 15674 9384 15674 0 _0039_
rlabel metal1 10166 20298 10166 20298 0 _0040_
rlabel metal2 8602 20094 8602 20094 0 _0041_
rlabel metal1 11178 21896 11178 21896 0 _0042_
rlabel metal2 9982 23256 9982 23256 0 _0043_
rlabel metal2 12282 24344 12282 24344 0 _0044_
rlabel metal1 13892 23834 13892 23834 0 _0045_
rlabel metal1 14122 25126 14122 25126 0 _0046_
rlabel metal2 12374 22440 12374 22440 0 _0047_
rlabel metal2 13662 21522 13662 21522 0 _0048_
rlabel metal1 13708 21658 13708 21658 0 _0049_
rlabel metal1 16146 14042 16146 14042 0 _0050_
rlabel metal2 15594 14178 15594 14178 0 _0051_
rlabel metal1 15088 12410 15088 12410 0 _0052_
rlabel metal1 2576 12614 2576 12614 0 _0053_
rlabel metal2 2438 10200 2438 10200 0 _0054_
rlabel metal2 2806 8092 2806 8092 0 _0055_
rlabel metal1 5382 5277 5382 5277 0 _0056_
rlabel metal2 5474 6120 5474 6120 0 _0057_
rlabel metal1 8464 10234 8464 10234 0 _0058_
rlabel metal2 10442 9758 10442 9758 0 _0059_
rlabel metal1 12519 3434 12519 3434 0 _0060_
rlabel metal2 14950 3230 14950 3230 0 _0061_
rlabel metal1 17940 4250 17940 4250 0 _0062_
rlabel metal2 18078 8670 18078 8670 0 _0063_
rlabel metal1 17342 3162 17342 3162 0 _0064_
rlabel metal1 18814 10744 18814 10744 0 _0065_
rlabel metal2 18446 10506 18446 10506 0 _0066_
rlabel metal1 13800 8058 13800 8058 0 _0067_
rlabel metal1 13156 2890 13156 2890 0 _0068_
rlabel metal2 13478 13124 13478 13124 0 _0069_
rlabel metal2 21390 13906 21390 13906 0 _0070_
rlabel metal2 21850 5848 21850 5848 0 _0071_
rlabel metal1 22349 3502 22349 3502 0 _0072_
rlabel metal2 20930 4318 20930 4318 0 _0073_
rlabel metal1 21075 8942 21075 8942 0 _0074_
rlabel metal1 21942 8296 21942 8296 0 _0075_
rlabel metal2 21482 6562 21482 6562 0 _0076_
rlabel metal1 21850 10744 21850 10744 0 _0077_
rlabel metal2 21482 12002 21482 12002 0 _0078_
rlabel metal2 21022 13736 21022 13736 0 _0079_
rlabel metal1 19734 22406 19734 22406 0 _0080_
rlabel metal2 21022 23086 21022 23086 0 _0081_
rlabel metal1 20976 24650 20976 24650 0 _0082_
rlabel metal1 8149 25194 8149 25194 0 _0083_
rlabel metal1 9016 25466 9016 25466 0 _0084_
rlabel metal2 11822 25432 11822 25432 0 _0085_
rlabel metal2 21482 25432 21482 25432 0 _0086_
rlabel metal1 22487 23766 22487 23766 0 _0087_
rlabel metal2 18814 25704 18814 25704 0 _0088_
rlabel metal1 10534 24378 10534 24378 0 _0089_
rlabel metal2 24426 19550 24426 19550 0 _0090_
rlabel metal2 24978 18462 24978 18462 0 _0091_
rlabel metal2 24518 13736 24518 13736 0 _0092_
rlabel metal2 23690 13022 23690 13022 0 _0093_
rlabel metal1 22540 15334 22540 15334 0 _0094_
rlabel metal1 24748 14586 24748 14586 0 _0095_
rlabel metal1 25208 16422 25208 16422 0 _0096_
rlabel metal2 24702 10812 24702 10812 0 _0097_
rlabel metal2 25346 8942 25346 8942 0 _0098_
rlabel metal2 23690 9758 23690 9758 0 _0099_
rlabel metal1 17480 13702 17480 13702 0 _0100_
rlabel metal1 19320 13158 19320 13158 0 _0101_
rlabel metal1 11260 16762 11260 16762 0 _0102_
rlabel metal1 4462 12274 4462 12274 0 _0103_
rlabel metal1 12834 15674 12834 15674 0 _0104_
rlabel metal1 10902 14008 10902 14008 0 _0105_
rlabel metal1 3312 19278 3312 19278 0 _0106_
rlabel metal1 3910 21488 3910 21488 0 _0107_
rlabel metal1 2201 22202 2201 22202 0 _0108_
rlabel metal1 2254 19482 2254 19482 0 _0109_
rlabel metal1 19596 18870 19596 18870 0 _0110_
rlabel metal1 20976 17306 20976 17306 0 _0111_
rlabel metal1 21298 20570 21298 20570 0 _0112_
rlabel metal1 21068 18666 21068 18666 0 _0113_
rlabel metal2 18078 19550 18078 19550 0 _0114_
rlabel metal1 11822 19720 11822 19720 0 _0115_
rlabel metal2 11822 18394 11822 18394 0 _0116_
rlabel metal1 10258 18394 10258 18394 0 _0117_
rlabel metal1 6118 14450 6118 14450 0 _0118_
rlabel metal2 3128 12036 3128 12036 0 _0119_
rlabel metal1 3082 12920 3082 12920 0 _0120_
rlabel metal1 7084 12954 7084 12954 0 _0121_
rlabel metal1 6709 3706 6709 3706 0 _0122_
rlabel metal1 8096 2958 8096 2958 0 _0123_
rlabel metal1 10120 4046 10120 4046 0 _0124_
rlabel metal1 5152 3162 5152 3162 0 _0125_
rlabel metal1 11500 5270 11500 5270 0 _0126_
rlabel metal1 11638 6426 11638 6426 0 _0127_
rlabel metal2 18354 6766 18354 6766 0 _0128_
rlabel metal1 14996 7786 14996 7786 0 _0129_
rlabel via1 9423 11322 9423 11322 0 _0130_
rlabel metal1 8924 13498 8924 13498 0 _0131_
rlabel metal1 12581 12342 12581 12342 0 _0132_
rlabel metal1 12328 13226 12328 13226 0 _0133_
rlabel metal1 9154 25194 9154 25194 0 _0134_
rlabel metal2 12006 25398 12006 25398 0 _0135_
rlabel metal2 20378 25670 20378 25670 0 _0136_
rlabel metal1 21666 24208 21666 24208 0 _0137_
rlabel metal1 18998 25296 18998 25296 0 _0138_
rlabel metal1 10626 24208 10626 24208 0 _0139_
rlabel metal1 23966 18802 23966 18802 0 _0140_
rlabel metal2 23966 18326 23966 18326 0 _0141_
rlabel metal2 24886 19380 24886 19380 0 _0142_
rlabel metal1 24656 17850 24656 17850 0 _0143_
rlabel metal1 24886 12954 24886 12954 0 _0144_
rlabel metal1 23920 12410 23920 12410 0 _0145_
rlabel metal1 23920 14586 23920 14586 0 _0146_
rlabel metal1 25162 14416 25162 14416 0 _0147_
rlabel metal1 25116 16558 25116 16558 0 _0148_
rlabel metal1 24886 11084 24886 11084 0 _0149_
rlabel metal1 25530 9588 25530 9588 0 _0150_
rlabel metal1 23552 10030 23552 10030 0 _0151_
rlabel metal2 17986 13430 17986 13430 0 _0152_
rlabel metal1 19274 12410 19274 12410 0 _0153_
rlabel metal1 16376 8398 16376 8398 0 _0154_
rlabel metal2 12558 13702 12558 13702 0 _0155_
rlabel metal1 12696 12206 12696 12206 0 _0156_
rlabel metal1 9338 13294 9338 13294 0 _0157_
rlabel metal1 9614 11798 9614 11798 0 _0158_
rlabel metal1 15272 8466 15272 8466 0 _0159_
rlabel metal2 12190 13209 12190 13209 0 _0160_
rlabel metal1 18400 6970 18400 6970 0 _0161_
rlabel metal1 11684 6290 11684 6290 0 _0162_
rlabel metal1 11316 4794 11316 4794 0 _0163_
rlabel metal1 5934 2992 5934 2992 0 _0164_
rlabel metal1 10442 3706 10442 3706 0 _0165_
rlabel metal1 8602 3706 8602 3706 0 _0166_
rlabel metal1 7682 3706 7682 3706 0 _0167_
rlabel metal1 7406 12852 7406 12852 0 _0168_
rlabel metal1 3128 13906 3128 13906 0 _0169_
rlabel metal1 3588 13294 3588 13294 0 _0170_
rlabel metal2 19918 18190 19918 18190 0 _0171_
rlabel metal1 6716 14994 6716 14994 0 _0172_
rlabel metal1 10626 18258 10626 18258 0 _0173_
rlabel metal2 12006 18938 12006 18938 0 _0174_
rlabel metal2 11454 20060 11454 20060 0 _0175_
rlabel metal1 18216 18938 18216 18938 0 _0176_
rlabel metal1 21758 18394 21758 18394 0 _0177_
rlabel metal1 21712 20434 21712 20434 0 _0178_
rlabel metal1 21574 17170 21574 17170 0 _0179_
rlabel metal1 19366 17850 19366 17850 0 _0180_
rlabel metal1 2622 19414 2622 19414 0 _0181_
rlabel metal1 21160 16014 21160 16014 0 _0182_
rlabel metal1 2691 22610 2691 22610 0 _0183_
rlabel metal2 3818 22440 3818 22440 0 _0184_
rlabel metal2 3818 19686 3818 19686 0 _0185_
rlabel metal1 11316 13906 11316 13906 0 _0186_
rlabel metal1 13156 15470 13156 15470 0 _0187_
rlabel metal1 5336 12410 5336 12410 0 _0188_
rlabel metal1 11454 17170 11454 17170 0 _0189_
rlabel metal1 14076 14586 14076 14586 0 _0190_
rlabel metal2 22034 15096 22034 15096 0 _0191_
rlabel metal1 14628 22542 14628 22542 0 _0192_
rlabel metal1 5520 19414 5520 19414 0 _0193_
rlabel metal1 2898 17238 2898 17238 0 _0194_
rlabel metal1 2990 16150 2990 16150 0 _0195_
rlabel metal2 3082 17782 3082 17782 0 _0196_
rlabel metal1 3956 16014 3956 16014 0 _0197_
rlabel metal1 4186 16116 4186 16116 0 _0198_
rlabel metal1 3588 15062 3588 15062 0 _0199_
rlabel metal2 2806 15232 2806 15232 0 _0200_
rlabel metal1 2438 14484 2438 14484 0 _0201_
rlabel metal2 8786 7684 8786 7684 0 _0202_
rlabel metal2 8556 7310 8556 7310 0 _0203_
rlabel metal1 7958 7990 7958 7990 0 _0204_
rlabel metal2 8694 7361 8694 7361 0 _0205_
rlabel metal1 8142 4726 8142 4726 0 _0206_
rlabel metal1 6854 6834 6854 6834 0 _0207_
rlabel metal2 7498 6290 7498 6290 0 _0208_
rlabel metal1 7498 6154 7498 6154 0 _0209_
rlabel metal2 8970 5916 8970 5916 0 _0210_
rlabel metal1 9154 7412 9154 7412 0 _0211_
rlabel metal1 9384 6970 9384 6970 0 _0212_
rlabel metal1 8970 6834 8970 6834 0 _0213_
rlabel metal1 8602 6732 8602 6732 0 _0214_
rlabel metal1 7590 7344 7590 7344 0 _0215_
rlabel metal2 4830 8092 4830 8092 0 _0216_
rlabel metal1 4140 9418 4140 9418 0 _0217_
rlabel metal1 5336 9010 5336 9010 0 _0218_
rlabel metal1 6992 10506 6992 10506 0 _0219_
rlabel metal1 6992 11254 6992 11254 0 _0220_
rlabel metal1 6578 11118 6578 11118 0 _0221_
rlabel metal1 5060 10642 5060 10642 0 _0222_
rlabel metal2 5382 10812 5382 10812 0 _0223_
rlabel metal1 5428 9486 5428 9486 0 _0224_
rlabel metal1 6256 7854 6256 7854 0 _0225_
rlabel metal2 8142 17952 8142 17952 0 _0226_
rlabel via1 8786 17647 8786 17647 0 _0227_
rlabel metal1 8004 17306 8004 17306 0 _0228_
rlabel metal1 7682 17680 7682 17680 0 _0229_
rlabel metal1 20700 16558 20700 16558 0 _0230_
rlabel metal1 21482 16524 21482 16524 0 _0231_
rlabel metal1 21850 16762 21850 16762 0 _0232_
rlabel metal1 16054 15640 16054 15640 0 _0233_
rlabel metal1 8234 17646 8234 17646 0 _0234_
rlabel metal1 8510 17680 8510 17680 0 _0235_
rlabel metal1 7268 19346 7268 19346 0 _0236_
rlabel metal2 6578 21692 6578 21692 0 _0237_
rlabel metal1 6486 19414 6486 19414 0 _0238_
rlabel metal2 6854 19550 6854 19550 0 _0239_
rlabel metal1 7544 19822 7544 19822 0 _0240_
rlabel metal1 5382 21522 5382 21522 0 _0241_
rlabel metal1 4692 22950 4692 22950 0 _0242_
rlabel metal1 5704 21998 5704 21998 0 _0243_
rlabel metal1 5796 21862 5796 21862 0 _0244_
rlabel metal1 7498 21556 7498 21556 0 _0245_
rlabel metal1 5980 21998 5980 21998 0 _0246_
rlabel metal1 7222 21522 7222 21522 0 _0247_
rlabel metal1 6693 22066 6693 22066 0 _0248_
rlabel metal1 5704 23086 5704 23086 0 _0249_
rlabel metal1 5658 22202 5658 22202 0 _0250_
rlabel metal2 5934 23324 5934 23324 0 _0251_
rlabel metal1 6946 21998 6946 21998 0 _0252_
rlabel metal1 8280 21862 8280 21862 0 _0253_
rlabel metal1 15640 17578 15640 17578 0 _0254_
rlabel metal2 15410 18496 15410 18496 0 _0255_
rlabel metal1 16836 19346 16836 19346 0 _0256_
rlabel metal1 14674 18938 14674 18938 0 _0257_
rlabel metal1 17112 18190 17112 18190 0 _0258_
rlabel metal1 15778 18224 15778 18224 0 _0259_
rlabel metal1 16974 18768 16974 18768 0 _0260_
rlabel metal1 16422 18666 16422 18666 0 _0261_
rlabel metal1 16330 19380 16330 19380 0 _0262_
rlabel metal1 17250 22576 17250 22576 0 _0263_
rlabel metal1 17296 21590 17296 21590 0 _0264_
rlabel metal1 17618 22746 17618 22746 0 _0265_
rlabel metal1 17020 22678 17020 22678 0 _0266_
rlabel metal1 17940 22542 17940 22542 0 _0267_
rlabel metal1 16284 24174 16284 24174 0 _0268_
rlabel metal1 17020 24174 17020 24174 0 _0269_
rlabel metal1 16928 23494 16928 23494 0 _0270_
rlabel metal1 17296 24922 17296 24922 0 _0271_
rlabel metal1 17158 24242 17158 24242 0 _0272_
rlabel metal1 16928 24786 16928 24786 0 _0273_
rlabel metal1 16008 20502 16008 20502 0 _0274_
rlabel metal1 16790 21522 16790 21522 0 _0275_
rlabel metal2 17066 22406 17066 22406 0 _0276_
rlabel metal1 17066 21658 17066 21658 0 _0277_
rlabel metal1 17158 20026 17158 20026 0 _0278_
rlabel metal1 15088 18734 15088 18734 0 _0279_
rlabel metal1 14858 18666 14858 18666 0 _0280_
rlabel metal2 15594 18054 15594 18054 0 _0281_
rlabel metal1 14950 18394 14950 18394 0 _0282_
rlabel metal2 14674 18853 14674 18853 0 _0283_
rlabel metal1 15732 19346 15732 19346 0 _0284_
rlabel metal2 15824 19210 15824 19210 0 _0285_
rlabel metal1 14352 19686 14352 19686 0 _0286_
rlabel metal1 5106 8908 5106 8908 0 _0287_
rlabel metal1 5474 9554 5474 9554 0 _0288_
rlabel metal1 3634 9894 3634 9894 0 _0289_
rlabel metal1 4600 8942 4600 8942 0 _0290_
rlabel metal1 6210 7344 6210 7344 0 _0291_
rlabel metal1 8142 6324 8142 6324 0 _0292_
rlabel metal1 7866 6426 7866 6426 0 _0293_
rlabel metal1 7636 6970 7636 6970 0 _0294_
rlabel metal1 14214 6188 14214 6188 0 _0295_
rlabel metal1 16514 6358 16514 6358 0 _0296_
rlabel metal1 17388 6154 17388 6154 0 _0297_
rlabel metal2 17158 5950 17158 5950 0 _0298_
rlabel metal1 19550 5746 19550 5746 0 _0299_
rlabel metal1 18538 5576 18538 5576 0 _0300_
rlabel metal1 18354 5678 18354 5678 0 _0301_
rlabel metal1 17434 5882 17434 5882 0 _0302_
rlabel metal2 16146 6460 16146 6460 0 _0303_
rlabel metal1 15088 4114 15088 4114 0 _0304_
rlabel metal1 13754 4080 13754 4080 0 _0305_
rlabel metal2 13754 4828 13754 4828 0 _0306_
rlabel metal1 15640 5746 15640 5746 0 _0307_
rlabel metal1 15824 4590 15824 4590 0 _0308_
rlabel metal2 15318 6086 15318 6086 0 _0309_
rlabel metal1 15226 4556 15226 4556 0 _0310_
rlabel metal2 15870 5066 15870 5066 0 _0311_
rlabel metal1 15042 6256 15042 6256 0 _0312_
rlabel metal1 14766 9554 14766 9554 0 _0313_
rlabel metal2 14766 10710 14766 10710 0 _0314_
rlabel metal1 14996 10166 14996 10166 0 _0315_
rlabel metal1 15594 9588 15594 9588 0 _0316_
rlabel metal1 15962 9520 15962 9520 0 _0317_
rlabel metal1 13478 9690 13478 9690 0 _0318_
rlabel metal1 12926 10744 12926 10744 0 _0319_
rlabel metal2 12098 10472 12098 10472 0 _0320_
rlabel metal1 13248 10098 13248 10098 0 _0321_
rlabel metal2 11914 9095 11914 9095 0 _0322_
rlabel metal1 12604 10030 12604 10030 0 _0323_
rlabel metal1 11638 9554 11638 9554 0 _0324_
rlabel metal1 15732 9554 15732 9554 0 _0325_
rlabel metal1 12834 10132 12834 10132 0 _0326_
rlabel metal1 12236 9554 12236 9554 0 _0327_
rlabel metal1 12880 9690 12880 9690 0 _0328_
rlabel metal2 4370 8670 4370 8670 0 _0329_
rlabel metal1 20838 16150 20838 16150 0 _0330_
rlabel metal1 19044 16694 19044 16694 0 _0331_
rlabel metal2 19182 16150 19182 16150 0 _0332_
rlabel metal1 21574 16422 21574 16422 0 _0333_
rlabel metal1 20470 16660 20470 16660 0 _0334_
rlabel metal1 19366 16728 19366 16728 0 _0335_
rlabel metal1 17158 16116 17158 16116 0 _0336_
rlabel metal1 14674 13872 14674 13872 0 _0337_
rlabel metal1 8602 19822 8602 19822 0 _0338_
rlabel metal2 8602 16796 8602 16796 0 _0339_
rlabel metal1 8326 16524 8326 16524 0 _0340_
rlabel metal1 7360 18326 7360 18326 0 _0341_
rlabel metal2 7682 18564 7682 18564 0 _0342_
rlabel metal1 8004 18122 8004 18122 0 _0343_
rlabel metal1 8326 19754 8326 19754 0 _0344_
rlabel metal1 9430 19788 9430 19788 0 _0345_
rlabel metal1 7314 19482 7314 19482 0 _0346_
rlabel via2 15134 19907 15134 19907 0 _0347_
rlabel metal1 7728 20026 7728 20026 0 _0348_
rlabel metal1 7314 21590 7314 21590 0 _0349_
rlabel metal1 7038 22202 7038 22202 0 _0350_
rlabel metal1 8004 22406 8004 22406 0 _0351_
rlabel metal1 8694 22066 8694 22066 0 _0352_
rlabel metal1 6210 21556 6210 21556 0 _0353_
rlabel metal1 7130 22746 7130 22746 0 _0354_
rlabel metal1 8142 22542 8142 22542 0 _0355_
rlabel metal1 8464 22610 8464 22610 0 _0356_
rlabel metal1 5888 21590 5888 21590 0 _0357_
rlabel metal1 7590 23698 7590 23698 0 _0358_
rlabel metal1 9890 23664 9890 23664 0 _0359_
rlabel metal2 15962 25126 15962 25126 0 _0360_
rlabel metal1 15778 23834 15778 23834 0 _0361_
rlabel metal1 14858 24140 14858 24140 0 _0362_
rlabel metal1 14582 24208 14582 24208 0 _0363_
rlabel metal1 16192 24718 16192 24718 0 _0364_
rlabel viali 15226 24172 15226 24172 0 _0365_
rlabel metal1 15456 24378 15456 24378 0 _0366_
rlabel metal2 16238 23290 16238 23290 0 _0367_
rlabel metal2 14214 22610 14214 22610 0 _0368_
rlabel metal1 13202 22746 13202 22746 0 _0369_
rlabel metal1 12374 23120 12374 23120 0 _0370_
rlabel metal1 17112 22950 17112 22950 0 _0371_
rlabel metal1 17480 22066 17480 22066 0 _0372_
rlabel metal1 17296 21930 17296 21930 0 _0373_
rlabel metal2 15962 22406 15962 22406 0 _0374_
rlabel metal1 14674 22746 14674 22746 0 _0375_
rlabel metal1 15778 19890 15778 19890 0 _0376_
rlabel metal1 14858 19788 14858 19788 0 _0377_
rlabel metal1 15778 19686 15778 19686 0 _0378_
rlabel metal1 14858 20026 14858 20026 0 _0379_
rlabel metal1 15962 17714 15962 17714 0 _0380_
rlabel metal1 15870 17612 15870 17612 0 _0381_
rlabel metal1 16606 17306 16606 17306 0 _0382_
rlabel metal1 15456 16966 15456 16966 0 _0383_
rlabel metal2 15778 16422 15778 16422 0 _0384_
rlabel metal1 15226 15470 15226 15470 0 _0385_
rlabel via1 15398 14994 15398 14994 0 _0386_
rlabel metal1 15134 17102 15134 17102 0 _0387_
rlabel metal1 14858 16626 14858 16626 0 _0388_
rlabel metal1 14996 14994 14996 14994 0 _0389_
rlabel metal2 14766 14416 14766 14416 0 _0390_
rlabel metal1 15456 12886 15456 12886 0 _0391_
rlabel metal1 6808 11322 6808 11322 0 _0392_
rlabel metal1 7544 11866 7544 11866 0 _0393_
rlabel metal1 7774 9996 7774 9996 0 _0394_
rlabel metal1 5566 10098 5566 10098 0 _0395_
rlabel metal2 5474 10676 5474 10676 0 _0396_
rlabel metal1 4738 10676 4738 10676 0 _0397_
rlabel metal1 4140 9486 4140 9486 0 _0398_
rlabel metal1 3910 9010 3910 9010 0 _0399_
rlabel metal1 1978 8500 1978 8500 0 _0400_
rlabel via1 3730 8466 3730 8466 0 _0401_
rlabel metal1 3726 7922 3726 7922 0 _0402_
rlabel metal1 4140 6766 4140 6766 0 _0403_
rlabel metal2 4692 6290 4692 6290 0 _0404_
rlabel metal1 6946 7718 6946 7718 0 _0405_
rlabel metal1 8096 6766 8096 6766 0 _0406_
rlabel metal1 6670 7310 6670 7310 0 _0407_
rlabel metal1 5842 6324 5842 6324 0 _0408_
rlabel metal2 7314 7956 7314 7956 0 _0409_
rlabel metal1 7820 8398 7820 8398 0 _0410_
rlabel metal1 7912 9690 7912 9690 0 _0411_
rlabel metal2 8326 7582 8326 7582 0 _0412_
rlabel metal1 9660 8058 9660 8058 0 _0413_
rlabel metal2 9338 8772 9338 8772 0 _0414_
rlabel metal1 9798 8806 9798 8806 0 _0415_
rlabel metal1 9292 6290 9292 6290 0 _0416_
rlabel metal2 9890 6732 9890 6732 0 _0417_
rlabel metal1 9430 6256 9430 6256 0 _0418_
rlabel metal1 9752 6222 9752 6222 0 _0419_
rlabel metal1 14996 5202 14996 5202 0 _0420_
rlabel metal1 15272 5202 15272 5202 0 _0421_
rlabel metal1 14030 5236 14030 5236 0 _0422_
rlabel metal1 14674 5134 14674 5134 0 _0423_
rlabel metal2 14766 4692 14766 4692 0 _0424_
rlabel metal1 16238 4658 16238 4658 0 _0425_
rlabel metal1 15962 5168 15962 5168 0 _0426_
rlabel metal1 17342 5644 17342 5644 0 _0427_
rlabel metal1 18032 6086 18032 6086 0 _0428_
rlabel metal2 18170 8330 18170 8330 0 _0429_
rlabel metal1 17434 8602 17434 8602 0 _0430_
rlabel metal1 16422 5780 16422 5780 0 _0431_
rlabel metal2 16514 5372 16514 5372 0 _0432_
rlabel metal1 16836 5270 16836 5270 0 _0433_
rlabel metal1 16376 9418 16376 9418 0 _0434_
rlabel metal1 15916 10030 15916 10030 0 _0435_
rlabel metal1 16008 10234 16008 10234 0 _0436_
rlabel metal1 16882 9962 16882 9962 0 _0437_
rlabel metal2 15410 10676 15410 10676 0 _0438_
rlabel metal1 15962 11186 15962 11186 0 _0439_
rlabel metal1 14030 9520 14030 9520 0 _0440_
rlabel metal1 13708 9894 13708 9894 0 _0441_
rlabel metal1 13248 8942 13248 8942 0 _0442_
rlabel metal1 12098 8500 12098 8500 0 _0443_
rlabel viali 11914 8468 11914 8468 0 _0444_
rlabel metal1 20792 14994 20792 14994 0 _0445_
rlabel metal1 21620 7378 21620 7378 0 _0446_
rlabel metal2 20930 3332 20930 3332 0 _0447_
rlabel metal1 19596 15062 19596 15062 0 _0448_
rlabel metal1 21942 3162 21942 3162 0 _0449_
rlabel metal1 19182 8942 19182 8942 0 _0450_
rlabel metal1 21482 8976 21482 8976 0 _0451_
rlabel metal1 20792 5338 20792 5338 0 _0452_
rlabel metal1 21298 11186 21298 11186 0 _0453_
rlabel metal1 21850 11832 21850 11832 0 _0454_
rlabel metal1 20148 13294 20148 13294 0 _0455_
rlabel metal2 18354 21692 18354 21692 0 _0456_
rlabel metal1 20700 21658 20700 21658 0 _0457_
rlabel metal2 20930 23460 20930 23460 0 _0458_
rlabel metal1 21206 25772 21206 25772 0 _0459_
rlabel metal2 6394 25092 6394 25092 0 _0460_
rlabel metal1 7820 24174 7820 24174 0 _0461_
rlabel metal1 9982 25466 9982 25466 0 _0462_
rlabel metal1 21666 24820 21666 24820 0 _0463_
rlabel metal1 21160 23834 21160 23834 0 _0464_
rlabel metal1 17848 25466 17848 25466 0 _0465_
rlabel metal1 8694 25262 8694 25262 0 _0466_
rlabel metal1 23736 20434 23736 20434 0 _0467_
rlabel metal1 23276 19346 23276 19346 0 _0468_
rlabel metal1 23598 17238 23598 17238 0 _0469_
rlabel metal1 22954 10234 22954 10234 0 _0470_
rlabel metal1 24196 15674 24196 15674 0 _0471_
rlabel metal2 21942 14688 21942 14688 0 _0472_
rlabel metal2 22862 16354 22862 16354 0 _0473_
rlabel metal1 24518 11118 24518 11118 0 _0474_
rlabel metal1 25438 8942 25438 8942 0 _0475_
rlabel metal1 23506 8874 23506 8874 0 _0476_
rlabel metal1 16514 12954 16514 12954 0 _0477_
rlabel metal1 18446 12274 18446 12274 0 _0478_
rlabel metal1 14398 17578 14398 17578 0 _0479_
rlabel metal2 13294 18666 13294 18666 0 _0480_
rlabel metal1 10764 17714 10764 17714 0 _0481_
rlabel metal1 12006 16218 12006 16218 0 _0482_
rlabel metal2 13754 14858 13754 14858 0 _0483_
rlabel metal1 12742 7514 12742 7514 0 _0484_
rlabel metal1 10810 11526 10810 11526 0 _0485_
rlabel metal1 10948 2890 10948 2890 0 _0486_
rlabel metal1 8786 12682 8786 12682 0 _0487_
rlabel metal2 11362 11968 11362 11968 0 _0488_
rlabel metal1 12006 20026 12006 20026 0 _0489_
rlabel metal2 10902 15844 10902 15844 0 _0490_
rlabel metal1 19826 12818 19826 12818 0 _0491_
rlabel via1 5566 16694 5566 16694 0 _0492_
rlabel metal1 5842 15130 5842 15130 0 _0493_
rlabel metal1 6072 16558 6072 16558 0 _0494_
rlabel metal1 6440 16558 6440 16558 0 _0495_
rlabel metal1 2438 17102 2438 17102 0 _0496_
rlabel metal1 3358 16218 3358 16218 0 _0497_
rlabel metal1 3128 14382 3128 14382 0 _0498_
rlabel metal2 12650 16796 12650 16796 0 _0499_
rlabel metal1 5152 13906 5152 13906 0 _0500_
rlabel metal1 12581 15470 12581 15470 0 _0501_
rlabel metal1 11730 14960 11730 14960 0 _0502_
rlabel metal1 18446 19890 18446 19890 0 _0503_
rlabel metal1 20194 19958 20194 19958 0 _0504_
rlabel metal1 3726 20400 3726 20400 0 _0505_
rlabel metal1 3404 20910 3404 20910 0 _0506_
rlabel metal1 2530 21114 2530 21114 0 _0507_
rlabel metal1 5382 19856 5382 19856 0 _0508_
rlabel metal1 19872 19822 19872 19822 0 _0509_
rlabel metal1 21252 18258 21252 18258 0 _0510_
rlabel metal1 21252 21114 21252 21114 0 _0511_
rlabel metal1 21850 19856 21850 19856 0 _0512_
rlabel metal1 19688 18734 19688 18734 0 _0513_
rlabel metal2 13018 20604 13018 20604 0 _0514_
rlabel metal1 10028 16014 10028 16014 0 _0515_
rlabel metal1 10488 15946 10488 15946 0 _0516_
rlabel metal1 10764 16762 10764 16762 0 _0517_
rlabel metal1 10626 16218 10626 16218 0 _0518_
rlabel metal1 6302 13906 6302 13906 0 _0519_
rlabel metal1 5106 11730 5106 11730 0 _0520_
rlabel metal1 5106 13294 5106 13294 0 _0521_
rlabel metal1 7130 13294 7130 13294 0 _0522_
rlabel metal1 7130 3026 7130 3026 0 _0523_
rlabel metal1 10672 3502 10672 3502 0 _0524_
rlabel metal1 10350 4624 10350 4624 0 _0525_
rlabel metal1 6118 3026 6118 3026 0 _0526_
rlabel metal1 17756 6766 17756 6766 0 _0527_
rlabel metal1 18676 13158 18676 13158 0 _0528_
rlabel metal1 11592 5678 11592 5678 0 _0529_
rlabel metal1 12489 6290 12489 6290 0 _0530_
rlabel metal1 18584 6902 18584 6902 0 _0531_
rlabel metal1 15778 7344 15778 7344 0 _0532_
rlabel metal1 10810 10234 10810 10234 0 _0533_
rlabel metal1 10580 14042 10580 14042 0 _0534_
rlabel metal1 12282 11696 12282 11696 0 _0535_
rlabel metal1 19366 14586 19366 14586 0 _0536_
rlabel metal1 18446 14960 18446 14960 0 _0537_
rlabel metal2 9982 15300 9982 15300 0 _0538_
rlabel metal2 12742 25024 12742 25024 0 _0539_
rlabel metal1 13294 22134 13294 22134 0 _0540_
rlabel metal1 10350 20434 10350 20434 0 _0541_
rlabel metal1 8786 20876 8786 20876 0 _0542_
rlabel metal1 10948 21658 10948 21658 0 _0543_
rlabel metal1 10212 22746 10212 22746 0 _0544_
rlabel metal2 12466 24310 12466 24310 0 _0545_
rlabel metal1 13892 23698 13892 23698 0 _0546_
rlabel metal2 13202 25092 13202 25092 0 _0547_
rlabel metal1 12489 21998 12489 21998 0 _0548_
rlabel metal2 13846 21386 13846 21386 0 _0549_
rlabel metal1 13340 21522 13340 21522 0 _0550_
rlabel metal1 1932 10574 1932 10574 0 _0551_
rlabel metal2 2438 7038 2438 7038 0 _0552_
rlabel metal1 15594 12954 15594 12954 0 _0553_
rlabel metal1 15640 13906 15640 13906 0 _0554_
rlabel metal1 14720 12206 14720 12206 0 _0555_
rlabel metal2 2438 12342 2438 12342 0 _0556_
rlabel metal1 2714 10608 2714 10608 0 _0557_
rlabel metal2 2530 7990 2530 7990 0 _0558_
rlabel viali 5198 6291 5198 6291 0 _0559_
rlabel viali 5658 6767 5658 6767 0 _0560_
rlabel metal1 8510 10030 8510 10030 0 _0561_
rlabel metal1 9752 9146 9752 9146 0 _0562_
rlabel metal1 13386 7922 13386 7922 0 _0563_
rlabel metal1 17066 2584 17066 2584 0 _0564_
rlabel metal1 12742 2482 12742 2482 0 _0565_
rlabel metal1 15088 2618 15088 2618 0 _0566_
rlabel metal1 18078 4080 18078 4080 0 _0567_
rlabel metal2 17986 8500 17986 8500 0 _0568_
rlabel metal1 17296 3026 17296 3026 0 _0569_
rlabel metal1 18952 10642 18952 10642 0 _0570_
rlabel metal1 18630 11152 18630 11152 0 _0571_
rlabel metal1 13938 7888 13938 7888 0 _0572_
rlabel metal1 13432 3026 13432 3026 0 _0573_
rlabel metal1 13570 12410 13570 12410 0 _0574_
rlabel metal1 20424 12750 20424 12750 0 _0575_
rlabel metal1 20516 12682 20516 12682 0 _0576_
rlabel metal1 21528 12954 21528 12954 0 _0577_
rlabel metal1 21298 5882 21298 5882 0 _0578_
rlabel metal1 22310 4182 22310 4182 0 _0579_
rlabel metal1 20930 4590 20930 4590 0 _0580_
rlabel metal2 20838 9078 20838 9078 0 _0581_
rlabel metal1 21758 8466 21758 8466 0 _0582_
rlabel metal1 21528 6290 21528 6290 0 _0583_
rlabel metal1 21436 10234 21436 10234 0 _0584_
rlabel metal1 21666 11696 21666 11696 0 _0585_
rlabel metal1 21068 12954 21068 12954 0 _0586_
rlabel metal1 18630 24174 18630 24174 0 _0587_
rlabel metal2 19550 23392 19550 23392 0 _0588_
rlabel metal1 19688 22610 19688 22610 0 _0589_
rlabel metal1 20562 23290 20562 23290 0 _0590_
rlabel metal1 20792 24378 20792 24378 0 _0591_
rlabel metal1 8510 25228 8510 25228 0 _0592_
rlabel metal1 8510 15062 8510 15062 0 clk
rlabel metal1 15686 20944 15686 20944 0 clknet_0_clk
rlabel metal1 2093 7922 2093 7922 0 clknet_3_0__leaf_clk
rlabel metal2 1426 11152 1426 11152 0 clknet_3_1__leaf_clk
rlabel metal1 15778 3468 15778 3468 0 clknet_3_2__leaf_clk
rlabel metal2 14122 13838 14122 13838 0 clknet_3_3__leaf_clk
rlabel metal1 2714 19414 2714 19414 0 clknet_3_4__leaf_clk
rlabel metal1 2438 21590 2438 21590 0 clknet_3_5__leaf_clk
rlabel metal1 16606 16014 16606 16014 0 clknet_3_6__leaf_clk
rlabel metal1 18262 21114 18262 21114 0 clknet_3_7__leaf_clk
rlabel metal2 4646 17918 4646 17918 0 cycle_reg.bit0.BitData
rlabel metal1 4186 17714 4186 17714 0 cycle_reg.bit0.BitOut
rlabel metal1 4646 18360 4646 18360 0 cycle_reg.bit1.BitData
rlabel metal1 4186 17612 4186 17612 0 cycle_reg.bit1.BitOut
rlabel metal1 2024 17714 2024 17714 0 cycle_reg.bit2.BitData
rlabel metal1 4002 17680 4002 17680 0 cycle_reg.bit2.BitOut
rlabel metal2 4278 16456 4278 16456 0 cycle_reg.bit3.BitData
rlabel metal1 3588 16626 3588 16626 0 cycle_reg.bit3.BitOut
rlabel metal1 2070 14586 2070 14586 0 cycle_reg.bit4.BitData
rlabel metal2 3358 15164 3358 15164 0 cycle_reg.bit4.BitOut
rlabel metal2 18722 1520 18722 1520 0 err
rlabel metal1 21574 15980 21574 15980 0 net1
rlabel metal2 18262 25874 18262 25874 0 net10
rlabel metal1 2530 2482 2530 2482 0 net100
rlabel metal1 17756 18258 17756 18258 0 net101
rlabel metal2 25254 22882 25254 22882 0 net102
rlabel metal1 22494 2346 22494 2346 0 net103
rlabel metal1 24610 25262 24610 25262 0 net104
rlabel metal3 15295 2652 15295 2652 0 net105
rlabel metal1 2300 13226 2300 13226 0 net106
rlabel metal1 1518 9520 1518 9520 0 net107
rlabel metal1 1518 3128 1518 3128 0 net108
rlabel metal1 7498 4556 7498 4556 0 net109
rlabel metal1 6900 26010 6900 26010 0 net11
rlabel metal2 2162 19890 2162 19890 0 net110
rlabel metal1 7452 7922 7452 7922 0 net111
rlabel metal2 10120 17238 10120 17238 0 net112
rlabel metal2 2622 19380 2622 19380 0 net113
rlabel metal2 5198 2210 5198 2210 0 net114
rlabel metal1 5474 1870 5474 1870 0 net115
rlabel metal1 20286 6698 20286 6698 0 net116
rlabel metal2 15088 17204 15088 17204 0 net117
rlabel metal2 17802 3026 17802 3026 0 net118
rlabel metal1 20654 12308 20654 12308 0 net119
rlabel metal2 22218 7718 22218 7718 0 net12
rlabel metal1 19872 5202 19872 5202 0 net120
rlabel metal1 4462 19346 4462 19346 0 net121
rlabel metal1 1518 8432 1518 8432 0 net122
rlabel metal1 5382 1836 5382 1836 0 net123
rlabel metal2 10166 20128 10166 20128 0 net124
rlabel metal1 2139 3434 2139 3434 0 net125
rlabel metal1 10902 21862 10902 21862 0 net126
rlabel metal2 9844 12716 9844 12716 0 net127
rlabel metal1 19366 24820 19366 24820 0 net128
rlabel metal2 16882 25874 16882 25874 0 net129
rlabel metal1 24886 21658 24886 21658 0 net13
rlabel metal1 2438 25806 2438 25806 0 net130
rlabel metal2 19366 2108 19366 2108 0 net131
rlabel metal2 19642 15436 19642 15436 0 net132
rlabel metal2 20654 16830 20654 16830 0 net133
rlabel metal1 4278 16422 4278 16422 0 net134
rlabel metal1 3266 15436 3266 15436 0 net135
rlabel metal1 5474 18870 5474 18870 0 net136
rlabel metal1 5934 18938 5934 18938 0 net137
rlabel metal1 17158 7514 17158 7514 0 net138
rlabel metal1 7498 20468 7498 20468 0 net139
rlabel metal2 2714 22797 2714 22797 0 net14
rlabel metal1 24564 8874 24564 8874 0 net140
rlabel metal1 14168 24174 14168 24174 0 net141
rlabel metal1 7820 8058 7820 8058 0 net142
rlabel metal1 4370 10642 4370 10642 0 net143
rlabel metal1 15410 24752 15410 24752 0 net144
rlabel metal1 12972 8942 12972 8942 0 net145
rlabel metal1 14306 4794 14306 4794 0 net146
rlabel metal1 10396 25194 10396 25194 0 net147
rlabel metal1 11638 17000 11638 17000 0 net148
rlabel metal1 7774 24684 7774 24684 0 net149
rlabel metal1 24426 17646 24426 17646 0 net15
rlabel metal1 9706 18258 9706 18258 0 net150
rlabel metal1 23368 16218 23368 16218 0 net151
rlabel metal1 22586 3094 22586 3094 0 net152
rlabel metal1 12466 12682 12466 12682 0 net153
rlabel metal1 22494 17306 22494 17306 0 net154
rlabel metal1 16284 8602 16284 8602 0 net155
rlabel metal1 18446 16422 18446 16422 0 net156
rlabel metal1 19872 16762 19872 16762 0 net157
rlabel metal1 19727 15674 19727 15674 0 net158
rlabel metal1 12466 4454 12466 4454 0 net159
rlabel metal2 12466 1972 12466 1972 0 net16
rlabel metal1 3956 22610 3956 22610 0 net160
rlabel metal1 21896 22950 21896 22950 0 net161
rlabel metal2 4554 6511 4554 6511 0 net162
rlabel metal1 4784 21862 4784 21862 0 net163
rlabel metal1 19320 6630 19320 6630 0 net164
rlabel metal2 22126 3774 22126 3774 0 net165
rlabel metal2 8418 3740 8418 3740 0 net166
rlabel metal1 25806 22406 25806 22406 0 net17
rlabel metal1 19481 2006 19481 2006 0 net18
rlabel metal2 1886 16541 1886 16541 0 net19
rlabel metal1 18308 21998 18308 21998 0 net2
rlabel metal1 25070 11322 25070 11322 0 net20
rlabel metal1 24978 3706 24978 3706 0 net21
rlabel metal1 25070 3638 25070 3638 0 net22
rlabel metal1 19274 2618 19274 2618 0 net23
rlabel metal1 16836 12886 16836 12886 0 net24
rlabel metal1 11270 2312 11270 2312 0 net25
rlabel metal1 23322 3162 23322 3162 0 net26
rlabel metal2 1472 18156 1472 18156 0 net27
rlabel metal2 22908 25670 22908 25670 0 net28
rlabel metal2 1610 4505 1610 4505 0 net29
rlabel metal1 22264 2550 22264 2550 0 net3
rlabel metal1 6578 11560 6578 11560 0 net30
rlabel metal2 25300 14484 25300 14484 0 net31
rlabel via2 20562 13243 20562 13243 0 net32
rlabel metal2 11914 17425 11914 17425 0 net33
rlabel metal1 23322 26214 23322 26214 0 net34
rlabel metal1 23598 17646 23598 17646 0 net35
rlabel metal2 18538 19006 18538 19006 0 net36
rlabel metal1 12558 20570 12558 20570 0 net37
rlabel metal2 13110 20009 13110 20009 0 net38
rlabel metal2 13018 19703 13018 19703 0 net39
rlabel metal2 21436 17204 21436 17204 0 net4
rlabel metal1 18170 26418 18170 26418 0 net40
rlabel metal1 1610 14280 1610 14280 0 net41
rlabel metal1 3404 14042 3404 14042 0 net42
rlabel metal1 22954 1938 22954 1938 0 net43
rlabel metal1 23230 17646 23230 17646 0 net44
rlabel metal1 9752 3026 9752 3026 0 net45
rlabel metal2 9338 3162 9338 3162 0 net46
rlabel metal1 12650 3536 12650 3536 0 net47
rlabel metal1 6762 2958 6762 2958 0 net48
rlabel metal2 5474 3570 5474 3570 0 net49
rlabel metal1 3772 7242 3772 7242 0 net5
rlabel metal1 12558 7446 12558 7446 0 net50
rlabel metal1 19642 2550 19642 2550 0 net51
rlabel metal1 25392 26350 25392 26350 0 net52
rlabel metal2 2162 15912 2162 15912 0 net53
rlabel metal1 14398 16490 14398 16490 0 net54
rlabel metal2 20010 2108 20010 2108 0 net55
rlabel via2 11914 12835 11914 12835 0 net56
rlabel metal2 11914 14314 11914 14314 0 net57
rlabel metal1 10166 12750 10166 12750 0 net58
rlabel metal1 4876 2618 4876 2618 0 net59
rlabel metal1 5290 5032 5290 5032 0 net6
rlabel metal1 17250 21012 17250 21012 0 net60
rlabel metal1 3910 19890 3910 19890 0 net61
rlabel metal1 4278 19822 4278 19822 0 net62
rlabel via2 1610 17051 1610 17051 0 net63
rlabel metal2 10718 13022 10718 13022 0 net64
rlabel metal1 1610 23732 1610 23732 0 net65
rlabel metal1 20424 20434 20424 20434 0 net66
rlabel metal2 14076 23732 14076 23732 0 net67
rlabel via2 1518 19363 1518 19363 0 net68
rlabel metal1 21896 23154 21896 23154 0 net69
rlabel metal1 9430 2550 9430 2550 0 net7
rlabel metal2 21114 24769 21114 24769 0 net70
rlabel metal2 8234 25874 8234 25874 0 net71
rlabel metal2 10258 26078 10258 26078 0 net72
rlabel metal1 2530 21352 2530 21352 0 net73
rlabel metal2 22218 24378 22218 24378 0 net74
rlabel metal1 23966 23494 23966 23494 0 net75
rlabel metal1 18814 25806 18814 25806 0 net76
rlabel metal2 2530 18972 2530 18972 0 net77
rlabel metal2 23138 3842 23138 3842 0 net78
rlabel metal1 25530 19482 25530 19482 0 net79
rlabel metal2 23046 26112 23046 26112 0 net8
rlabel metal1 19642 6392 19642 6392 0 net80
rlabel metal1 23322 10166 23322 10166 0 net81
rlabel metal1 1656 26282 1656 26282 0 net82
rlabel metal1 1886 16082 1886 16082 0 net83
rlabel metal1 24932 15130 24932 15130 0 net84
rlabel metal1 25668 25194 25668 25194 0 net85
rlabel metal2 2162 10523 2162 10523 0 net86
rlabel metal1 25392 8330 25392 8330 0 net87
rlabel metal1 22080 9384 22080 9384 0 net88
rlabel metal1 25024 2414 25024 2414 0 net89
rlabel via2 1610 23579 1610 23579 0 net9
rlabel metal1 17480 13498 17480 13498 0 net90
rlabel metal1 21942 2448 21942 2448 0 net91
rlabel via2 3910 2363 3910 2363 0 net92
rlabel via2 1518 10659 1518 10659 0 net93
rlabel metal2 23046 4352 23046 4352 0 net94
rlabel metal2 21942 10608 21942 10608 0 net95
rlabel via2 2070 3043 2070 3043 0 net96
rlabel metal1 21528 2414 21528 2414 0 net97
rlabel via2 1518 18275 1518 18275 0 net98
rlabel metal1 24150 7446 24150 7446 0 net99
rlabel metal3 820 7548 820 7548 0 ok
rlabel metal1 19274 16082 19274 16082 0 reg32_denom.bit0.BitOut
rlabel metal1 22080 17510 22080 17510 0 reg32_denom.bit1.BitOut
rlabel metal2 17434 21114 17434 21114 0 reg32_denom.bit10.BitOut
rlabel metal2 22310 18496 22310 18496 0 reg32_denom.bit11.BitOut
rlabel metal1 18630 18802 18630 18802 0 reg32_denom.bit12.BitOut
rlabel metal1 12926 20026 12926 20026 0 reg32_denom.bit13.BitOut
rlabel metal1 13064 18394 13064 18394 0 reg32_denom.bit14.BitOut
rlabel metal2 11638 19074 11638 19074 0 reg32_denom.bit15.BitOut
rlabel metal2 7314 14586 7314 14586 0 reg32_denom.bit16.BitOut
rlabel metal1 4416 13158 4416 13158 0 reg32_denom.bit17.BitOut
rlabel metal1 4508 12954 4508 12954 0 reg32_denom.bit18.BitOut
rlabel metal1 5934 12070 5934 12070 0 reg32_denom.bit19.BitOut
rlabel metal2 8418 13498 8418 13498 0 reg32_denom.bit2.BitOut
rlabel metal1 7866 4590 7866 4590 0 reg32_denom.bit20.BitOut
rlabel metal1 8418 5848 8418 5848 0 reg32_denom.bit21.BitOut
rlabel metal1 10166 6936 10166 6936 0 reg32_denom.bit22.BitOut
rlabel metal2 6808 2958 6808 2958 0 reg32_denom.bit23.BitOut
rlabel metal2 13294 4828 13294 4828 0 reg32_denom.bit24.BitOut
rlabel metal1 12834 6970 12834 6970 0 reg32_denom.bit25.BitOut
rlabel via1 19826 6834 19826 6834 0 reg32_denom.bit26.BitOut
rlabel metal1 16330 8058 16330 8058 0 reg32_denom.bit27.BitOut
rlabel metal1 10488 11322 10488 11322 0 reg32_denom.bit28.BitOut
rlabel metal1 13938 16422 13938 16422 0 reg32_denom.bit29.BitOut
rlabel metal2 9062 18258 9062 18258 0 reg32_denom.bit3.BitOut
rlabel metal1 12052 12750 12052 12750 0 reg32_denom.bit30.BitOut
rlabel metal1 12190 14042 12190 14042 0 reg32_denom.bit31.BitOut
rlabel metal1 4462 19244 4462 19244 0 reg32_denom.bit4.BitOut
rlabel metal2 5198 21182 5198 21182 0 reg32_denom.bit5.BitOut
rlabel metal1 3726 22542 3726 22542 0 reg32_denom.bit6.BitOut
rlabel metal1 4646 19686 4646 19686 0 reg32_denom.bit7.BitOut
rlabel metal1 20654 19482 20654 19482 0 reg32_denom.bit8.BitOut
rlabel metal1 15272 13498 15272 13498 0 reg32_denom.bit9.BitOut
rlabel metal2 20746 14620 20746 14620 0 reg32_result.bit0.BitData
rlabel metal2 21206 6460 21206 6460 0 reg32_result.bit1.BitData
rlabel metal1 19090 21658 19090 21658 0 reg32_result.bit10.BitData
rlabel metal1 20930 22202 20930 22202 0 reg32_result.bit11.BitData
rlabel metal1 19918 23834 19918 23834 0 reg32_result.bit12.BitData
rlabel metal1 6486 25194 6486 25194 0 reg32_result.bit13.BitData
rlabel metal1 8418 24378 8418 24378 0 reg32_result.bit14.BitData
rlabel metal1 11316 25330 11316 25330 0 reg32_result.bit15.BitData
rlabel metal1 21252 24922 21252 24922 0 reg32_result.bit16.BitData
rlabel metal2 22034 23936 22034 23936 0 reg32_result.bit17.BitData
rlabel metal1 18170 25976 18170 25976 0 reg32_result.bit18.BitData
rlabel metal1 8878 24854 8878 24854 0 reg32_result.bit19.BitData
rlabel metal1 21298 3400 21298 3400 0 reg32_result.bit2.BitData
rlabel metal1 23736 19414 23736 19414 0 reg32_result.bit20.BitData
rlabel metal1 23414 18360 23414 18360 0 reg32_result.bit21.BitData
rlabel metal2 24058 15470 24058 15470 0 reg32_result.bit22.BitData
rlabel metal1 22908 11322 22908 11322 0 reg32_result.bit23.BitData
rlabel metal1 22632 15402 22632 15402 0 reg32_result.bit24.BitData
rlabel metal1 22954 14586 22954 14586 0 reg32_result.bit25.BitData
rlabel metal1 23920 16150 23920 16150 0 reg32_result.bit26.BitData
rlabel metal1 23598 10744 23598 10744 0 reg32_result.bit27.BitData
rlabel metal1 24058 8568 24058 8568 0 reg32_result.bit28.BitData
rlabel metal1 23138 9146 23138 9146 0 reg32_result.bit29.BitData
rlabel metal1 21022 4046 21022 4046 0 reg32_result.bit3.BitData
rlabel metal1 16422 13226 16422 13226 0 reg32_result.bit30.BitData
rlabel metal1 18308 12410 18308 12410 0 reg32_result.bit31.BitData
rlabel metal1 19310 9146 19310 9146 0 reg32_result.bit4.BitData
rlabel metal1 21160 7922 21160 7922 0 reg32_result.bit5.BitData
rlabel metal1 20746 6426 20746 6426 0 reg32_result.bit6.BitData
rlabel metal1 20102 10744 20102 10744 0 reg32_result.bit7.BitData
rlabel metal1 20562 12138 20562 12138 0 reg32_result.bit8.BitData
rlabel metal1 19964 13498 19964 13498 0 reg32_result.bit9.BitData
rlabel metal1 19688 16082 19688 16082 0 reg32_work.bit0.BitData
rlabel metal1 17434 16014 17434 16014 0 reg32_work.bit1.BitData
rlabel metal1 11914 22712 11914 22712 0 reg32_work.bit10.BitData
rlabel metal1 14250 22202 14250 22202 0 reg32_work.bit11.BitData
rlabel metal1 14214 20842 14214 20842 0 reg32_work.bit12.BitData
rlabel metal1 16192 15402 16192 15402 0 reg32_work.bit13.BitData
rlabel metal1 15180 14450 15180 14450 0 reg32_work.bit14.BitData
rlabel metal1 14352 13226 14352 13226 0 reg32_work.bit15.BitData
rlabel metal1 1702 12104 1702 12104 0 reg32_work.bit16.BitData
rlabel metal1 2231 10098 2231 10098 0 reg32_work.bit17.BitData
rlabel metal1 1840 7786 1840 7786 0 reg32_work.bit18.BitData
rlabel metal1 4462 5134 4462 5134 0 reg32_work.bit19.BitData
rlabel metal1 8050 16150 8050 16150 0 reg32_work.bit2.BitData
rlabel metal1 5244 5746 5244 5746 0 reg32_work.bit20.BitData
rlabel metal1 7682 10234 7682 10234 0 reg32_work.bit21.BitData
rlabel metal1 9200 9622 9200 9622 0 reg32_work.bit22.BitData
rlabel metal1 11355 3706 11355 3706 0 reg32_work.bit23.BitData
rlabel metal1 14168 3094 14168 3094 0 reg32_work.bit24.BitData
rlabel metal1 16376 4522 16376 4522 0 reg32_work.bit25.BitData
rlabel metal2 17526 8602 17526 8602 0 reg32_work.bit26.BitData
rlabel metal1 16100 3434 16100 3434 0 reg32_work.bit27.BitData
rlabel metal1 16376 10574 16376 10574 0 reg32_work.bit28.BitData
rlabel metal1 17112 10098 17112 10098 0 reg32_work.bit29.BitData
rlabel metal1 8694 20026 8694 20026 0 reg32_work.bit3.BitData
rlabel metal2 12742 8670 12742 8670 0 reg32_work.bit30.BitData
rlabel metal2 11822 4964 11822 4964 0 reg32_work.bit31.BitData
rlabel metal1 7590 19414 7590 19414 0 reg32_work.bit4.BitData
rlabel metal1 8832 21930 8832 21930 0 reg32_work.bit5.BitData
rlabel metal1 8832 22746 8832 22746 0 reg32_work.bit6.BitData
rlabel metal1 9545 23834 9545 23834 0 reg32_work.bit7.BitData
rlabel metal1 13846 24378 13846 24378 0 reg32_work.bit8.BitData
rlabel metal1 14766 24922 14766 24922 0 reg32_work.bit9.BitData
rlabel metal3 820 23868 820 23868 0 reset
rlabel metal1 24978 13260 24978 13260 0 start
rlabel metal1 5014 15402 5014 15402 0 u1.d
rlabel metal1 16790 14484 16790 14484 0 u1.q
<< properties >>
string FIXED_BBOX 0 0 27037 29181
<< end >>
