// This is the unpowered netlist.
module divider (clk,
    err,
    ok,
    reset,
    start,
    A,
    B,
    D,
    R);
 input clk;
 output err;
 output ok;
 input reset;
 input start;
 input [31:0] A;
 input [31:0] B;
 output [31:0] D;
 output [31:0] R;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire \cycle_reg.bit0.BitData ;
 wire \cycle_reg.bit0.BitOut ;
 wire \cycle_reg.bit1.BitData ;
 wire \cycle_reg.bit1.BitOut ;
 wire \cycle_reg.bit2.BitData ;
 wire \cycle_reg.bit2.BitOut ;
 wire \cycle_reg.bit3.BitData ;
 wire \cycle_reg.bit3.BitOut ;
 wire \cycle_reg.bit4.BitData ;
 wire \cycle_reg.bit4.BitOut ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \reg32_denom.bit0.BitOut ;
 wire \reg32_denom.bit1.BitOut ;
 wire \reg32_denom.bit10.BitOut ;
 wire \reg32_denom.bit11.BitOut ;
 wire \reg32_denom.bit12.BitOut ;
 wire \reg32_denom.bit13.BitOut ;
 wire \reg32_denom.bit14.BitOut ;
 wire \reg32_denom.bit15.BitOut ;
 wire \reg32_denom.bit16.BitOut ;
 wire \reg32_denom.bit17.BitOut ;
 wire \reg32_denom.bit18.BitOut ;
 wire \reg32_denom.bit19.BitOut ;
 wire \reg32_denom.bit2.BitOut ;
 wire \reg32_denom.bit20.BitOut ;
 wire \reg32_denom.bit21.BitOut ;
 wire \reg32_denom.bit22.BitOut ;
 wire \reg32_denom.bit23.BitOut ;
 wire \reg32_denom.bit24.BitOut ;
 wire \reg32_denom.bit25.BitOut ;
 wire \reg32_denom.bit26.BitOut ;
 wire \reg32_denom.bit27.BitOut ;
 wire \reg32_denom.bit28.BitOut ;
 wire \reg32_denom.bit29.BitOut ;
 wire \reg32_denom.bit3.BitOut ;
 wire \reg32_denom.bit30.BitOut ;
 wire \reg32_denom.bit31.BitOut ;
 wire \reg32_denom.bit4.BitOut ;
 wire \reg32_denom.bit5.BitOut ;
 wire \reg32_denom.bit6.BitOut ;
 wire \reg32_denom.bit7.BitOut ;
 wire \reg32_denom.bit8.BitOut ;
 wire \reg32_denom.bit9.BitOut ;
 wire \reg32_result.bit0.BitData ;
 wire \reg32_result.bit1.BitData ;
 wire \reg32_result.bit10.BitData ;
 wire \reg32_result.bit11.BitData ;
 wire \reg32_result.bit12.BitData ;
 wire \reg32_result.bit13.BitData ;
 wire \reg32_result.bit14.BitData ;
 wire \reg32_result.bit15.BitData ;
 wire \reg32_result.bit16.BitData ;
 wire \reg32_result.bit17.BitData ;
 wire \reg32_result.bit18.BitData ;
 wire \reg32_result.bit19.BitData ;
 wire \reg32_result.bit2.BitData ;
 wire \reg32_result.bit20.BitData ;
 wire \reg32_result.bit21.BitData ;
 wire \reg32_result.bit22.BitData ;
 wire \reg32_result.bit23.BitData ;
 wire \reg32_result.bit24.BitData ;
 wire \reg32_result.bit25.BitData ;
 wire \reg32_result.bit26.BitData ;
 wire \reg32_result.bit27.BitData ;
 wire \reg32_result.bit28.BitData ;
 wire \reg32_result.bit29.BitData ;
 wire \reg32_result.bit3.BitData ;
 wire \reg32_result.bit30.BitData ;
 wire \reg32_result.bit31.BitData ;
 wire \reg32_result.bit4.BitData ;
 wire \reg32_result.bit5.BitData ;
 wire \reg32_result.bit6.BitData ;
 wire \reg32_result.bit7.BitData ;
 wire \reg32_result.bit8.BitData ;
 wire \reg32_result.bit9.BitData ;
 wire \reg32_work.bit0.BitData ;
 wire \reg32_work.bit1.BitData ;
 wire \reg32_work.bit10.BitData ;
 wire \reg32_work.bit11.BitData ;
 wire \reg32_work.bit12.BitData ;
 wire \reg32_work.bit13.BitData ;
 wire \reg32_work.bit14.BitData ;
 wire \reg32_work.bit15.BitData ;
 wire \reg32_work.bit16.BitData ;
 wire \reg32_work.bit17.BitData ;
 wire \reg32_work.bit18.BitData ;
 wire \reg32_work.bit19.BitData ;
 wire \reg32_work.bit2.BitData ;
 wire \reg32_work.bit20.BitData ;
 wire \reg32_work.bit21.BitData ;
 wire \reg32_work.bit22.BitData ;
 wire \reg32_work.bit23.BitData ;
 wire \reg32_work.bit24.BitData ;
 wire \reg32_work.bit25.BitData ;
 wire \reg32_work.bit26.BitData ;
 wire \reg32_work.bit27.BitData ;
 wire \reg32_work.bit28.BitData ;
 wire \reg32_work.bit29.BitData ;
 wire \reg32_work.bit3.BitData ;
 wire \reg32_work.bit30.BitData ;
 wire \reg32_work.bit31.BitData ;
 wire \reg32_work.bit4.BitData ;
 wire \reg32_work.bit5.BitData ;
 wire \reg32_work.bit6.BitData ;
 wire \reg32_work.bit7.BitData ;
 wire \reg32_work.bit8.BitData ;
 wire \reg32_work.bit9.BitData ;
 wire \u1.d ;
 wire \u1.q ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net83));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_96 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__clkbuf_4 _0593_ (.A(\u1.q ),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net64),
    .A1(\reg32_denom.bit9.BitOut ),
    .S(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0155_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net56),
    .A1(\reg32_denom.bit30.BitOut ),
    .S(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0156_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net58),
    .A1(\reg32_denom.bit3.BitOut ),
    .S(_0154_),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0599_ (.A(_0157_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net53),
    .A1(\reg32_denom.bit28.BitOut ),
    .S(_0154_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0601_ (.A(_0158_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net52),
    .A1(net155),
    .S(_0154_),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(_0159_),
    .X(_0129_));
 sky130_fd_sc_hd__buf_4 _0604_ (.A(\u1.q ),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(net51),
    .A1(net164),
    .S(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _0606_ (.A(_0161_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(net50),
    .A1(\reg32_denom.bit25.BitOut ),
    .S(_0160_),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(_0162_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0609_ (.A0(net49),
    .A1(net159),
    .S(_0160_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _0610_ (.A(_0163_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0611_ (.A0(net48),
    .A1(\reg32_denom.bit23.BitOut ),
    .S(_0160_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0164_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0613_ (.A0(net47),
    .A1(\reg32_denom.bit22.BitOut ),
    .S(_0160_),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(_0165_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0615_ (.A0(net46),
    .A1(\reg32_denom.bit21.BitOut ),
    .S(_0160_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0166_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0617_ (.A0(net45),
    .A1(net166),
    .S(_0160_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(_0167_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(net55),
    .A1(\reg32_denom.bit2.BitOut ),
    .S(_0160_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(_0168_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(net42),
    .A1(\reg32_denom.bit18.BitOut ),
    .S(_0160_),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0169_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(net41),
    .A1(\reg32_denom.bit17.BitOut ),
    .S(_0160_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0170_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_4 _0625_ (.A(\u1.q ),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(net40),
    .A1(\reg32_denom.bit16.BitOut ),
    .S(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0627_ (.A(_0172_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(net39),
    .A1(\reg32_denom.bit15.BitOut ),
    .S(_0171_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0629_ (.A(_0173_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(net38),
    .A1(\reg32_denom.bit14.BitOut ),
    .S(_0171_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0174_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(net37),
    .A1(\reg32_denom.bit13.BitOut ),
    .S(_0171_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _0633_ (.A(_0175_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(net36),
    .A1(\reg32_denom.bit12.BitOut ),
    .S(_0171_),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(_0176_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net35),
    .A1(\reg32_denom.bit11.BitOut ),
    .S(_0171_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _0637_ (.A(_0177_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(net34),
    .A1(\reg32_denom.bit10.BitOut ),
    .S(_0171_),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _0639_ (.A(_0178_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0640_ (.A0(net44),
    .A1(net154),
    .S(_0171_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0641_ (.A(_0179_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(net63),
    .A1(\reg32_denom.bit8.BitOut ),
    .S(_0171_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _0643_ (.A(_0180_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0644_ (.A0(net62),
    .A1(\reg32_denom.bit7.BitOut ),
    .S(_0171_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0645_ (.A(_0181_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_4 _0646_ (.A(\u1.q ),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(net61),
    .A1(net160),
    .S(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0183_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(net60),
    .A1(net163),
    .S(_0182_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0184_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0651_ (.A0(net59),
    .A1(\reg32_denom.bit4.BitOut ),
    .S(_0182_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _0652_ (.A(_0185_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0653_ (.A0(net57),
    .A1(\reg32_denom.bit31.BitOut ),
    .S(_0182_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0186_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(net54),
    .A1(\reg32_denom.bit29.BitOut ),
    .S(_0182_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _0656_ (.A(_0187_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0657_ (.A0(net43),
    .A1(\reg32_denom.bit19.BitOut ),
    .S(_0182_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(_0188_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(net33),
    .A1(\reg32_denom.bit0.BitOut ),
    .S(_0182_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0189_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _0661_ (.A(_0154_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_1 _0662_ (.A(_0190_),
    .B(net136),
    .Y(\cycle_reg.bit0.BitData ));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(\u1.q ),
    .Y(net132));
 sky130_fd_sc_hd__clkbuf_4 _0664_ (.A(\u1.q ),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_4 _0665_ (.A(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__o21ai_1 _0666_ (.A1(\cycle_reg.bit0.BitOut ),
    .A2(\cycle_reg.bit1.BitOut ),
    .B1(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__a21o_1 _0667_ (.A1(net136),
    .A2(net137),
    .B1(_0193_),
    .X(\cycle_reg.bit1.BitData ));
 sky130_fd_sc_hd__o21a_1 _0668_ (.A1(\cycle_reg.bit0.BitOut ),
    .A2(\cycle_reg.bit1.BitOut ),
    .B1(\cycle_reg.bit2.BitOut ),
    .X(_0194_));
 sky130_fd_sc_hd__or3_1 _0669_ (.A(\cycle_reg.bit0.BitOut ),
    .B(\cycle_reg.bit1.BitOut ),
    .C(\cycle_reg.bit2.BitOut ),
    .X(_0195_));
 sky130_fd_sc_hd__or3b_1 _0670_ (.A(_0194_),
    .B(net132),
    .C_N(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0671_ (.A(_0196_),
    .X(\cycle_reg.bit2.BitData ));
 sky130_fd_sc_hd__or2_1 _0672_ (.A(net134),
    .B(_0195_),
    .X(_0197_));
 sky130_fd_sc_hd__a21oi_1 _0673_ (.A1(net134),
    .A2(_0195_),
    .B1(net132),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(_0197_),
    .B(_0198_),
    .Y(\cycle_reg.bit3.BitData ));
 sky130_fd_sc_hd__nor2_1 _0675_ (.A(net135),
    .B(_0197_),
    .Y(_0199_));
 sky130_fd_sc_hd__a21o_1 _0676_ (.A1(\cycle_reg.bit4.BitOut ),
    .A2(_0197_),
    .B1(net132),
    .X(_0200_));
 sky130_fd_sc_hd__or2_1 _0677_ (.A(_0199_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0201_),
    .X(\cycle_reg.bit4.BitData ));
 sky130_fd_sc_hd__and2b_1 _0679_ (.A_N(net111),
    .B(\reg32_denom.bit21.BitOut ),
    .X(_0202_));
 sky130_fd_sc_hd__or2b_1 _0680_ (.A(\reg32_denom.bit21.BitOut ),
    .B_N(net111),
    .X(_0203_));
 sky130_fd_sc_hd__or2b_1 _0681_ (.A(_0202_),
    .B_N(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__or2b_2 _0682_ (.A(\reg32_denom.bit20.BitOut ),
    .B_N(net109),
    .X(_0205_));
 sky130_fd_sc_hd__or2b_1 _0683_ (.A(net109),
    .B_N(\reg32_denom.bit20.BitOut ),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _0684_ (.A(_0205_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__and2b_1 _0685_ (.A_N(net113),
    .B(\reg32_denom.bit23.BitOut ),
    .X(_0208_));
 sky130_fd_sc_hd__or2b_1 _0686_ (.A(\reg32_denom.bit23.BitOut ),
    .B_N(net113),
    .X(_0209_));
 sky130_fd_sc_hd__and2b_1 _0687_ (.A_N(_0208_),
    .B(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__and2b_1 _0689_ (.A_N(net112),
    .B(\reg32_denom.bit22.BitOut ),
    .X(_0212_));
 sky130_fd_sc_hd__or2b_1 _0690_ (.A(\reg32_denom.bit22.BitOut ),
    .B_N(net112),
    .X(_0213_));
 sky130_fd_sc_hd__or2b_1 _0691_ (.A(_0212_),
    .B_N(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__or4_1 _0692_ (.A(_0204_),
    .B(_0207_),
    .C(_0211_),
    .D(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__xor2_1 _0693_ (.A(\reg32_denom.bit19.BitOut ),
    .B(net108),
    .X(_0216_));
 sky130_fd_sc_hd__xnor2_1 _0694_ (.A(\reg32_denom.bit18.BitOut ),
    .B(net107),
    .Y(_0217_));
 sky130_fd_sc_hd__or2b_1 _0695_ (.A(_0216_),
    .B_N(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__or2b_1 _0696_ (.A(\reg32_denom.bit16.BitOut ),
    .B_N(net105),
    .X(_0219_));
 sky130_fd_sc_hd__or2b_1 _0697_ (.A(net105),
    .B_N(\reg32_denom.bit16.BitOut ),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _0698_ (.A(_0219_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__or2b_1 _0699_ (.A(net106),
    .B_N(\reg32_denom.bit17.BitOut ),
    .X(_0222_));
 sky130_fd_sc_hd__or2b_1 _0700_ (.A(\reg32_denom.bit17.BitOut ),
    .B_N(net106),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _0701_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__or3_1 _0702_ (.A(_0218_),
    .B(_0221_),
    .C(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__and2b_1 _0703_ (.A_N(net121),
    .B(\reg32_denom.bit3.BitOut ),
    .X(_0226_));
 sky130_fd_sc_hd__or2b_1 _0704_ (.A(\reg32_denom.bit2.BitOut ),
    .B_N(net110),
    .X(_0227_));
 sky130_fd_sc_hd__or2b_1 _0705_ (.A(net110),
    .B_N(\reg32_denom.bit2.BitOut ),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_1 _0706_ (.A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__or2b_1 _0707_ (.A(net91),
    .B_N(\reg32_denom.bit0.BitOut ),
    .X(_0230_));
 sky130_fd_sc_hd__or2b_1 _0708_ (.A(net99),
    .B_N(\reg32_denom.bit1.BitOut ),
    .X(_0231_));
 sky130_fd_sc_hd__and2b_1 _0709_ (.A_N(\reg32_denom.bit1.BitOut ),
    .B(net99),
    .X(_0232_));
 sky130_fd_sc_hd__a21oi_2 _0710_ (.A1(_0230_),
    .A2(_0231_),
    .B1(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__or3b_1 _0711_ (.A(\reg32_denom.bit2.BitOut ),
    .B(_0226_),
    .C_N(net110),
    .X(_0234_));
 sky130_fd_sc_hd__or2b_1 _0712_ (.A(\reg32_denom.bit3.BitOut ),
    .B_N(net121),
    .X(_0235_));
 sky130_fd_sc_hd__o311ai_2 _0713_ (.A1(_0226_),
    .A2(_0229_),
    .A3(_0233_),
    .B1(_0234_),
    .C1(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__and2b_1 _0714_ (.A_N(\reg32_denom.bit4.BitOut ),
    .B(net124),
    .X(_0237_));
 sky130_fd_sc_hd__and2b_1 _0715_ (.A_N(net124),
    .B(\reg32_denom.bit4.BitOut ),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_1 _0716_ (.A(_0237_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(_0236_),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__and2b_1 _0718_ (.A_N(\reg32_denom.bit6.BitOut ),
    .B(net126),
    .X(_0241_));
 sky130_fd_sc_hd__and2b_1 _0719_ (.A_N(net126),
    .B(\reg32_denom.bit6.BitOut ),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_1 _0720_ (.A(_0241_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_2 _0721_ (.A(\reg32_denom.bit7.BitOut ),
    .B(net127),
    .Y(_0244_));
 sky130_fd_sc_hd__or2b_1 _0722_ (.A(net125),
    .B_N(\reg32_denom.bit5.BitOut ),
    .X(_0245_));
 sky130_fd_sc_hd__and2b_1 _0723_ (.A_N(\reg32_denom.bit5.BitOut ),
    .B(net125),
    .X(_0246_));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__and4_1 _0725_ (.A(_0243_),
    .B(_0244_),
    .C(_0245_),
    .D(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(\reg32_denom.bit7.BitOut ),
    .Y(_0249_));
 sky130_fd_sc_hd__o2111a_1 _0727_ (.A1(_0237_),
    .A2(_0246_),
    .B1(_0245_),
    .C1(_0244_),
    .D1(_0243_),
    .X(_0250_));
 sky130_fd_sc_hd__o21a_1 _0728_ (.A1(_0249_),
    .A2(net127),
    .B1(_0241_),
    .X(_0251_));
 sky130_fd_sc_hd__a211o_1 _0729_ (.A1(_0249_),
    .A2(net127),
    .B1(_0250_),
    .C1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__a21oi_2 _0730_ (.A1(_0240_),
    .A2(_0248_),
    .B1(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__xor2_2 _0731_ (.A(\reg32_denom.bit14.BitOut ),
    .B(net103),
    .X(_0254_));
 sky130_fd_sc_hd__xor2_2 _0732_ (.A(\reg32_denom.bit15.BitOut ),
    .B(net104),
    .X(_0255_));
 sky130_fd_sc_hd__or2b_1 _0733_ (.A(net102),
    .B_N(\reg32_denom.bit13.BitOut ),
    .X(_0256_));
 sky130_fd_sc_hd__or2b_1 _0734_ (.A(\reg32_denom.bit13.BitOut ),
    .B_N(net102),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _0735_ (.A(_0256_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nor2b_1 _0736_ (.A(\reg32_denom.bit12.BitOut ),
    .B_N(net101),
    .Y(_0259_));
 sky130_fd_sc_hd__and2b_1 _0737_ (.A_N(net101),
    .B(\reg32_denom.bit12.BitOut ),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _0738_ (.A(_0259_),
    .B(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__or4_1 _0739_ (.A(_0254_),
    .B(_0255_),
    .C(_0258_),
    .D(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__xor2_1 _0740_ (.A(\reg32_denom.bit11.BitOut ),
    .B(net100),
    .X(_0263_));
 sky130_fd_sc_hd__and2b_1 _0741_ (.A_N(\reg32_denom.bit10.BitOut ),
    .B(net130),
    .X(_0264_));
 sky130_fd_sc_hd__and2b_1 _0742_ (.A_N(net130),
    .B(\reg32_denom.bit10.BitOut ),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _0743_ (.A(_0264_),
    .B(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _0744_ (.A(_0263_),
    .B(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__and2b_1 _0745_ (.A_N(\reg32_denom.bit8.BitOut ),
    .B(net128),
    .X(_0268_));
 sky130_fd_sc_hd__and2b_1 _0746_ (.A_N(net128),
    .B(\reg32_denom.bit8.BitOut ),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(_0268_),
    .B(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__and2b_1 _0748_ (.A_N(\reg32_denom.bit9.BitOut ),
    .B(net129),
    .X(_0271_));
 sky130_fd_sc_hd__or2b_1 _0749_ (.A(net129),
    .B_N(\reg32_denom.bit9.BitOut ),
    .X(_0272_));
 sky130_fd_sc_hd__or2b_1 _0750_ (.A(_0271_),
    .B_N(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__or3_1 _0751_ (.A(_0267_),
    .B(_0270_),
    .C(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(net100),
    .Y(_0275_));
 sky130_fd_sc_hd__o21ai_1 _0753_ (.A1(_0268_),
    .A2(_0271_),
    .B1(_0272_),
    .Y(_0276_));
 sky130_fd_sc_hd__a21bo_1 _0754_ (.A1(\reg32_denom.bit11.BitOut ),
    .A2(_0275_),
    .B1_N(_0264_),
    .X(_0277_));
 sky130_fd_sc_hd__o221a_1 _0755_ (.A1(\reg32_denom.bit11.BitOut ),
    .A2(_0275_),
    .B1(_0267_),
    .B2(_0276_),
    .C1(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(net104),
    .Y(_0279_));
 sky130_fd_sc_hd__a21bo_1 _0757_ (.A1(\reg32_denom.bit15.BitOut ),
    .A2(_0279_),
    .B1_N(net103),
    .X(_0280_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(_0257_),
    .Y(_0281_));
 sky130_fd_sc_hd__nor2_1 _0759_ (.A(_0254_),
    .B(_0255_),
    .Y(_0282_));
 sky130_fd_sc_hd__o211ai_1 _0760_ (.A1(_0281_),
    .A2(_0259_),
    .B1(_0282_),
    .C1(_0256_),
    .Y(_0283_));
 sky130_fd_sc_hd__o221a_1 _0761_ (.A1(\reg32_denom.bit15.BitOut ),
    .A2(_0279_),
    .B1(_0280_),
    .B2(\reg32_denom.bit14.BitOut ),
    .C1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__o21a_1 _0762_ (.A1(_0262_),
    .A2(_0278_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__o31a_2 _0763_ (.A1(_0253_),
    .A2(_0262_),
    .A3(_0274_),
    .B1(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(net108),
    .Y(_0287_));
 sky130_fd_sc_hd__a21bo_1 _0765_ (.A1(_0223_),
    .A2(_0219_),
    .B1_N(_0222_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(net107),
    .Y(_0289_));
 sky130_fd_sc_hd__a211o_1 _0767_ (.A1(\reg32_denom.bit19.BitOut ),
    .A2(_0287_),
    .B1(_0289_),
    .C1(\reg32_denom.bit18.BitOut ),
    .X(_0290_));
 sky130_fd_sc_hd__o221a_1 _0768_ (.A1(\reg32_denom.bit19.BitOut ),
    .A2(_0287_),
    .B1(_0288_),
    .B2(_0218_),
    .C1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _0769_ (.A(_0291_),
    .B(_0207_),
    .X(_0292_));
 sky130_fd_sc_hd__a311o_1 _0770_ (.A1(_0205_),
    .A2(_0203_),
    .A3(_0292_),
    .B1(_0202_),
    .C1(_0212_),
    .X(_0293_));
 sky130_fd_sc_hd__a31o_1 _0771_ (.A1(_0293_),
    .A2(_0213_),
    .A3(_0209_),
    .B1(_0208_),
    .X(_0294_));
 sky130_fd_sc_hd__o31ai_2 _0772_ (.A1(_0215_),
    .A2(_0225_),
    .A3(_0286_),
    .B1(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__and2b_1 _0773_ (.A_N(\reg32_denom.bit27.BitOut ),
    .B(net117),
    .X(_0296_));
 sky130_fd_sc_hd__or2b_1 _0774_ (.A(net117),
    .B_N(\reg32_denom.bit27.BitOut ),
    .X(_0297_));
 sky130_fd_sc_hd__and2b_1 _0775_ (.A_N(_0296_),
    .B(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__and2b_1 _0776_ (.A_N(\reg32_denom.bit26.BitOut ),
    .B(net116),
    .X(_0299_));
 sky130_fd_sc_hd__and2b_1 _0777_ (.A_N(net116),
    .B(\reg32_denom.bit26.BitOut ),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(_0299_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__and2_1 _0780_ (.A(_0298_),
    .B(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__and2b_1 _0781_ (.A_N(\reg32_denom.bit24.BitOut ),
    .B(net114),
    .X(_0304_));
 sky130_fd_sc_hd__and2b_1 _0782_ (.A_N(net114),
    .B(\reg32_denom.bit24.BitOut ),
    .X(_0305_));
 sky130_fd_sc_hd__nor2_1 _0783_ (.A(_0304_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__or2b_1 _0784_ (.A(\reg32_denom.bit25.BitOut ),
    .B_N(net115),
    .X(_0307_));
 sky130_fd_sc_hd__or2b_1 _0785_ (.A(net115),
    .B_N(\reg32_denom.bit25.BitOut ),
    .X(_0308_));
 sky130_fd_sc_hd__and4_1 _0786_ (.A(_0303_),
    .B(_0306_),
    .C(_0307_),
    .D(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__and2b_1 _0787_ (.A_N(\reg32_denom.bit25.BitOut ),
    .B(net115),
    .X(_0310_));
 sky130_fd_sc_hd__o21a_1 _0788_ (.A1(_0304_),
    .A2(_0310_),
    .B1(_0308_),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _0789_ (.A1(_0297_),
    .A2(_0299_),
    .B1(_0303_),
    .B2(_0311_),
    .C1(_0296_),
    .X(_0312_));
 sky130_fd_sc_hd__a21o_1 _0790_ (.A1(_0295_),
    .A2(_0309_),
    .B1(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__and2b_1 _0791_ (.A_N(net119),
    .B(\reg32_denom.bit29.BitOut ),
    .X(_0314_));
 sky130_fd_sc_hd__or2b_1 _0792_ (.A(\reg32_denom.bit29.BitOut ),
    .B_N(net119),
    .X(_0315_));
 sky130_fd_sc_hd__and2b_1 _0793_ (.A_N(_0314_),
    .B(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__xnor2_2 _0794_ (.A(\reg32_denom.bit28.BitOut ),
    .B(net118),
    .Y(_0317_));
 sky130_fd_sc_hd__nand3_2 _0795_ (.A(_0313_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__and2b_1 _0796_ (.A_N(\reg32_denom.bit30.BitOut ),
    .B(net120),
    .X(_0319_));
 sky130_fd_sc_hd__and2b_1 _0797_ (.A_N(net120),
    .B(\reg32_denom.bit30.BitOut ),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _0798_ (.A(_0319_),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__xor2_1 _0799_ (.A(\reg32_denom.bit31.BitOut ),
    .B(net122),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _0800_ (.A(_0321_),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(net122),
    .Y(_0324_));
 sky130_fd_sc_hd__or2b_1 _0802_ (.A(\reg32_denom.bit28.BitOut ),
    .B_N(net118),
    .X(_0325_));
 sky130_fd_sc_hd__a21o_1 _0803_ (.A1(_0315_),
    .A2(_0325_),
    .B1(_0314_),
    .X(_0326_));
 sky130_fd_sc_hd__a21bo_1 _0804_ (.A1(\reg32_denom.bit31.BitOut ),
    .A2(_0324_),
    .B1_N(_0319_),
    .X(_0327_));
 sky130_fd_sc_hd__o221a_1 _0805_ (.A1(\reg32_denom.bit31.BitOut ),
    .A2(_0324_),
    .B1(_0323_),
    .B2(_0326_),
    .C1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__o21ai_2 _0806_ (.A1(_0318_),
    .A2(_0323_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_4 _0807_ (.A(net133),
    .X(_0330_));
 sky130_fd_sc_hd__a21oi_1 _0808_ (.A1(net156),
    .A2(_0330_),
    .B1(net91),
    .Y(_0331_));
 sky130_fd_sc_hd__a31o_1 _0809_ (.A1(\reg32_denom.bit0.BitOut ),
    .A2(net91),
    .A3(_0330_),
    .B1(net132),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _0810_ (.A(net157),
    .B(_0332_),
    .Y(\reg32_work.bit0.BitData ));
 sky130_fd_sc_hd__or2b_1 _0811_ (.A(_0232_),
    .B_N(_0231_),
    .X(_0333_));
 sky130_fd_sc_hd__xnor2_1 _0812_ (.A(_0230_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(net99),
    .A1(_0334_),
    .S(net133),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _0814_ (.A(_0192_),
    .B(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _0815_ (.A(_0336_),
    .X(\reg32_work.bit1.BitData ));
 sky130_fd_sc_hd__clkbuf_4 _0816_ (.A(_0330_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_4 _0817_ (.A(_0330_),
    .X(_0338_));
 sky130_fd_sc_hd__xnor2_1 _0818_ (.A(_0229_),
    .B(_0233_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _0819_ (.A(_0338_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__o211a_1 _0820_ (.A1(net148),
    .A2(_0337_),
    .B1(_0340_),
    .C1(_0190_),
    .X(\reg32_work.bit2.BitData ));
 sky130_fd_sc_hd__o21ai_1 _0821_ (.A1(_0229_),
    .A2(_0233_),
    .B1(_0227_),
    .Y(_0341_));
 sky130_fd_sc_hd__and2b_1 _0822_ (.A_N(\reg32_denom.bit3.BitOut ),
    .B(net121),
    .X(_0342_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(_0342_),
    .B(_0226_),
    .Y(_0343_));
 sky130_fd_sc_hd__xnor2_1 _0824_ (.A(_0341_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(_0338_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__o211a_1 _0826_ (.A1(net150),
    .A2(_0337_),
    .B1(_0345_),
    .C1(_0190_),
    .X(\reg32_work.bit3.BitData ));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(_0236_),
    .B(_0239_),
    .Y(_0346_));
 sky130_fd_sc_hd__clkbuf_4 _0828_ (.A(net133),
    .X(_0347_));
 sky130_fd_sc_hd__o21ai_1 _0829_ (.A1(_0240_),
    .A2(_0346_),
    .B1(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__o211a_1 _0830_ (.A1(net139),
    .A2(_0337_),
    .B1(_0348_),
    .C1(_0190_),
    .X(\reg32_work.bit4.BitData ));
 sky130_fd_sc_hd__nand2_1 _0831_ (.A(_0245_),
    .B(_0247_),
    .Y(_0349_));
 sky130_fd_sc_hd__nor2_1 _0832_ (.A(_0237_),
    .B(_0240_),
    .Y(_0350_));
 sky130_fd_sc_hd__xnor2_1 _0833_ (.A(_0349_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(_0338_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__o211a_1 _0835_ (.A1(net125),
    .A2(_0337_),
    .B1(_0352_),
    .C1(_0190_),
    .X(\reg32_work.bit5.BitData ));
 sky130_fd_sc_hd__o31a_1 _0836_ (.A1(_0237_),
    .A2(_0240_),
    .A3(_0246_),
    .B1(_0245_),
    .X(_0353_));
 sky130_fd_sc_hd__xor2_1 _0837_ (.A(_0243_),
    .B(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(net126),
    .A1(_0354_),
    .S(net133),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _0839_ (.A(_0192_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(_0356_),
    .X(\reg32_work.bit6.BitData ));
 sky130_fd_sc_hd__a21o_1 _0841_ (.A1(_0243_),
    .A2(_0353_),
    .B1(_0241_),
    .X(_0357_));
 sky130_fd_sc_hd__xnor2_1 _0842_ (.A(_0244_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _0843_ (.A(_0338_),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__o211a_1 _0844_ (.A1(net127),
    .A2(_0337_),
    .B1(_0359_),
    .C1(_0190_),
    .X(\reg32_work.bit7.BitData ));
 sky130_fd_sc_hd__nor2_1 _0845_ (.A(_0253_),
    .B(_0270_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _0846_ (.A(_0253_),
    .B(_0270_),
    .Y(_0361_));
 sky130_fd_sc_hd__or2b_1 _0847_ (.A(_0360_),
    .B_N(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _0848_ (.A(_0338_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__o211a_1 _0849_ (.A1(net141),
    .A2(_0337_),
    .B1(_0363_),
    .C1(_0190_),
    .X(\reg32_work.bit8.BitData ));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(_0268_),
    .B(_0360_),
    .Y(_0364_));
 sky130_fd_sc_hd__xnor2_1 _0851_ (.A(_0273_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _0852_ (.A(_0338_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__o211a_1 _0853_ (.A1(net144),
    .A2(_0337_),
    .B1(_0366_),
    .C1(_0190_),
    .X(\reg32_work.bit9.BitData ));
 sky130_fd_sc_hd__o31a_1 _0854_ (.A1(_0268_),
    .A2(_0271_),
    .A3(_0360_),
    .B1(_0272_),
    .X(_0367_));
 sky130_fd_sc_hd__xnor2_1 _0855_ (.A(_0266_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(net130),
    .A1(_0368_),
    .S(net133),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _0857_ (.A(_0192_),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0858_ (.A(_0370_),
    .X(\reg32_work.bit10.BitData ));
 sky130_fd_sc_hd__inv_2 _0859_ (.A(_0266_),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_1 _0860_ (.A1(_0371_),
    .A2(_0367_),
    .B1(_0264_),
    .X(_0372_));
 sky130_fd_sc_hd__xnor2_1 _0861_ (.A(_0263_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(net100),
    .A1(_0373_),
    .S(net133),
    .X(_0374_));
 sky130_fd_sc_hd__and2_1 _0863_ (.A(_0192_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0864_ (.A(_0375_),
    .X(\reg32_work.bit11.BitData ));
 sky130_fd_sc_hd__or2_1 _0865_ (.A(_0253_),
    .B(_0274_),
    .X(_0376_));
 sky130_fd_sc_hd__and3_1 _0866_ (.A(_0261_),
    .B(_0278_),
    .C(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__a21oi_2 _0867_ (.A1(_0278_),
    .A2(_0376_),
    .B1(_0261_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_1 _0868_ (.A1(_0377_),
    .A2(_0378_),
    .B1(_0347_),
    .Y(_0379_));
 sky130_fd_sc_hd__o211a_1 _0869_ (.A1(net101),
    .A2(_0337_),
    .B1(_0379_),
    .C1(_0190_),
    .X(\reg32_work.bit12.BitData ));
 sky130_fd_sc_hd__o21ai_1 _0870_ (.A1(_0259_),
    .A2(_0378_),
    .B1(_0258_),
    .Y(_0380_));
 sky130_fd_sc_hd__or3_1 _0871_ (.A(_0258_),
    .B(_0259_),
    .C(_0378_),
    .X(_0381_));
 sky130_fd_sc_hd__o21ai_1 _0872_ (.A1(net102),
    .A2(_0330_),
    .B1(_0192_),
    .Y(_0382_));
 sky130_fd_sc_hd__a31oi_1 _0873_ (.A1(_0338_),
    .A2(_0380_),
    .A3(_0381_),
    .B1(_0382_),
    .Y(\reg32_work.bit13.BitData ));
 sky130_fd_sc_hd__o31ai_2 _0874_ (.A1(_0281_),
    .A2(_0259_),
    .A3(_0378_),
    .B1(_0256_),
    .Y(_0383_));
 sky130_fd_sc_hd__xor2_1 _0875_ (.A(_0254_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _0876_ (.A0(net103),
    .A1(_0384_),
    .S(net133),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0192_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _0878_ (.A(_0386_),
    .X(\reg32_work.bit14.BitData ));
 sky130_fd_sc_hd__or2b_1 _0879_ (.A(\reg32_denom.bit14.BitOut ),
    .B_N(net103),
    .X(_0387_));
 sky130_fd_sc_hd__o21a_1 _0880_ (.A1(_0254_),
    .A2(_0383_),
    .B1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0881_ (.A(_0255_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(_0338_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__clkbuf_4 _0883_ (.A(_0154_),
    .X(_0391_));
 sky130_fd_sc_hd__o211a_1 _0884_ (.A1(net104),
    .A2(_0337_),
    .B1(_0390_),
    .C1(_0391_),
    .X(\reg32_work.bit15.BitData ));
 sky130_fd_sc_hd__xnor2_1 _0885_ (.A(_0221_),
    .B(_0286_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0338_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__o211a_1 _0887_ (.A1(net153),
    .A2(_0337_),
    .B1(_0393_),
    .C1(_0391_),
    .X(\reg32_work.bit16.BitData ));
 sky130_fd_sc_hd__clkbuf_4 _0888_ (.A(_0330_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _0889_ (.A1(_0221_),
    .A2(_0286_),
    .B1(_0219_),
    .Y(_0395_));
 sky130_fd_sc_hd__xor2_1 _0890_ (.A(_0224_),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _0891_ (.A(_0347_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o211a_1 _0892_ (.A1(net143),
    .A2(_0394_),
    .B1(_0397_),
    .C1(_0391_),
    .X(\reg32_work.bit17.BitData ));
 sky130_fd_sc_hd__o31a_1 _0893_ (.A1(_0221_),
    .A2(_0224_),
    .A3(_0286_),
    .B1(_0288_),
    .X(_0398_));
 sky130_fd_sc_hd__xor2_1 _0894_ (.A(_0217_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _0895_ (.A0(_0289_),
    .A1(_0399_),
    .S(_0329_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(net132),
    .B(_0400_),
    .Y(\reg32_work.bit18.BitData ));
 sky130_fd_sc_hd__and2b_1 _0897_ (.A_N(_0398_),
    .B(_0217_),
    .X(_0401_));
 sky130_fd_sc_hd__o21ba_1 _0898_ (.A1(\reg32_denom.bit18.BitOut ),
    .A2(_0289_),
    .B1_N(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__xnor2_1 _0899_ (.A(_0216_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _0900_ (.A(_0347_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__o211a_1 _0901_ (.A1(net162),
    .A2(_0394_),
    .B1(_0404_),
    .C1(_0391_),
    .X(\reg32_work.bit19.BitData ));
 sky130_fd_sc_hd__or2_1 _0902_ (.A(_0225_),
    .B(_0286_),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _0903_ (.A1(_0291_),
    .A2(_0405_),
    .B1(_0207_),
    .X(_0406_));
 sky130_fd_sc_hd__nand3_1 _0904_ (.A(_0291_),
    .B(_0207_),
    .C(_0405_),
    .Y(_0407_));
 sky130_fd_sc_hd__a21bo_1 _0905_ (.A1(_0406_),
    .A2(_0407_),
    .B1_N(_0330_),
    .X(_0408_));
 sky130_fd_sc_hd__o211a_1 _0906_ (.A1(net109),
    .A2(_0394_),
    .B1(_0408_),
    .C1(_0391_),
    .X(\reg32_work.bit20.BitData ));
 sky130_fd_sc_hd__nand2_1 _0907_ (.A(_0205_),
    .B(_0406_),
    .Y(_0409_));
 sky130_fd_sc_hd__xor2_1 _0908_ (.A(_0204_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _0909_ (.A(_0347_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__o211a_1 _0910_ (.A1(net142),
    .A2(_0394_),
    .B1(_0411_),
    .C1(_0391_),
    .X(\reg32_work.bit21.BitData ));
 sky130_fd_sc_hd__a31o_1 _0911_ (.A1(_0205_),
    .A2(_0203_),
    .A3(_0406_),
    .B1(_0202_),
    .X(_0412_));
 sky130_fd_sc_hd__xor2_1 _0912_ (.A(_0214_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _0913_ (.A0(net112),
    .A1(_0413_),
    .S(_0329_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _0914_ (.A(_0154_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0415_),
    .X(\reg32_work.bit22.BitData ));
 sky130_fd_sc_hd__a311o_1 _0916_ (.A1(_0205_),
    .A2(_0203_),
    .A3(_0406_),
    .B1(_0214_),
    .C1(_0202_),
    .X(_0416_));
 sky130_fd_sc_hd__and3_1 _0917_ (.A(_0213_),
    .B(_0210_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a21o_1 _0918_ (.A1(_0213_),
    .A2(_0416_),
    .B1(_0210_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _0919_ (.A(_0347_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__o221a_1 _0920_ (.A1(net113),
    .A2(_0394_),
    .B1(_0417_),
    .B2(_0419_),
    .C1(_0192_),
    .X(\reg32_work.bit23.BitData ));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(_0295_),
    .B(_0306_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _0922_ (.A(_0295_),
    .B(_0306_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21ai_1 _0923_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0347_),
    .Y(_0422_));
 sky130_fd_sc_hd__o211a_1 _0924_ (.A1(net146),
    .A2(_0394_),
    .B1(_0422_),
    .C1(_0391_),
    .X(\reg32_work.bit24.BitData ));
 sky130_fd_sc_hd__nand2_1 _0925_ (.A(_0307_),
    .B(_0308_),
    .Y(_0423_));
 sky130_fd_sc_hd__nor2_1 _0926_ (.A(_0304_),
    .B(_0420_),
    .Y(_0424_));
 sky130_fd_sc_hd__xnor2_1 _0927_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(_0347_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__o211a_1 _0929_ (.A1(net115),
    .A2(_0394_),
    .B1(_0426_),
    .C1(_0391_),
    .X(\reg32_work.bit25.BitData ));
 sky130_fd_sc_hd__a31o_1 _0930_ (.A1(_0307_),
    .A2(_0308_),
    .A3(_0420_),
    .B1(_0311_),
    .X(_0427_));
 sky130_fd_sc_hd__xnor2_1 _0931_ (.A(_0301_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net116),
    .A1(_0428_),
    .S(net133),
    .X(_0429_));
 sky130_fd_sc_hd__and2_1 _0933_ (.A(_0154_),
    .B(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _0934_ (.A(_0430_),
    .X(\reg32_work.bit26.BitData ));
 sky130_fd_sc_hd__a21o_1 _0935_ (.A1(_0302_),
    .A2(_0427_),
    .B1(_0299_),
    .X(_0431_));
 sky130_fd_sc_hd__xnor2_1 _0936_ (.A(_0298_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__o21ai_1 _0937_ (.A1(net117),
    .A2(_0330_),
    .B1(_0192_),
    .Y(_0433_));
 sky130_fd_sc_hd__a21oi_1 _0938_ (.A1(_0394_),
    .A2(_0432_),
    .B1(_0433_),
    .Y(\reg32_work.bit27.BitData ));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(_0313_),
    .B(_0317_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _0940_ (.A(_0313_),
    .B(_0317_),
    .X(_0435_));
 sky130_fd_sc_hd__a21bo_1 _0941_ (.A1(_0434_),
    .A2(_0435_),
    .B1_N(_0330_),
    .X(_0436_));
 sky130_fd_sc_hd__o211a_1 _0942_ (.A1(net138),
    .A2(_0394_),
    .B1(_0436_),
    .C1(_0391_),
    .X(\reg32_work.bit28.BitData ));
 sky130_fd_sc_hd__and3_1 _0943_ (.A(_0316_),
    .B(_0325_),
    .C(_0434_),
    .X(_0437_));
 sky130_fd_sc_hd__a21o_1 _0944_ (.A1(_0325_),
    .A2(_0434_),
    .B1(_0316_),
    .X(_0438_));
 sky130_fd_sc_hd__nand2_1 _0945_ (.A(_0347_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__o221a_1 _0946_ (.A1(net119),
    .A2(_0338_),
    .B1(_0437_),
    .B2(_0439_),
    .C1(_0192_),
    .X(\reg32_work.bit29.BitData ));
 sky130_fd_sc_hd__and3_1 _0947_ (.A(_0318_),
    .B(_0321_),
    .C(_0326_),
    .X(_0440_));
 sky130_fd_sc_hd__a21oi_2 _0948_ (.A1(_0318_),
    .A2(_0326_),
    .B1(_0321_),
    .Y(_0441_));
 sky130_fd_sc_hd__o21ai_1 _0949_ (.A1(_0440_),
    .A2(_0441_),
    .B1(_0347_),
    .Y(_0442_));
 sky130_fd_sc_hd__o211a_1 _0950_ (.A1(net145),
    .A2(_0394_),
    .B1(_0442_),
    .C1(_0391_),
    .X(\reg32_work.bit30.BitData ));
 sky130_fd_sc_hd__nor2_1 _0951_ (.A(_0319_),
    .B(_0441_),
    .Y(_0443_));
 sky130_fd_sc_hd__o311a_1 _0952_ (.A1(\reg32_denom.bit31.BitOut ),
    .A2(_0319_),
    .A3(_0441_),
    .B1(net122),
    .C1(_0154_),
    .X(_0444_));
 sky130_fd_sc_hd__o21a_1 _0953_ (.A1(_0322_),
    .A2(_0443_),
    .B1(_0444_),
    .X(\reg32_work.bit31.BitData ));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net1),
    .A1(_0330_),
    .S(_0182_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0445_),
    .X(\reg32_result.bit0.BitData ));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net12),
    .A1(net67),
    .S(_0182_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0446_),
    .X(\reg32_result.bit1.BitData ));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(net23),
    .A1(net165),
    .S(_0182_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0447_),
    .X(\reg32_result.bit2.BitData ));
 sky130_fd_sc_hd__buf_4 _0960_ (.A(\u1.q ),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(net26),
    .A1(net152),
    .S(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _0962_ (.A(_0449_),
    .X(\reg32_result.bit3.BitData ));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(net27),
    .A1(net92),
    .S(_0448_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0450_),
    .X(\reg32_result.bit4.BitData ));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(net28),
    .A1(net93),
    .S(_0448_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(_0451_),
    .X(\reg32_result.bit5.BitData ));
 sky130_fd_sc_hd__mux2_1 _0967_ (.A0(net29),
    .A1(net94),
    .S(_0448_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0968_ (.A(_0452_),
    .X(\reg32_result.bit6.BitData ));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(net30),
    .A1(net95),
    .S(_0448_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0970_ (.A(_0453_),
    .X(\reg32_result.bit7.BitData ));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(net31),
    .A1(net96),
    .S(_0448_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0972_ (.A(_0454_),
    .X(\reg32_result.bit8.BitData ));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(net32),
    .A1(net97),
    .S(_0448_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(_0455_),
    .X(\reg32_result.bit9.BitData ));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(net2),
    .A1(net98),
    .S(_0448_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(_0456_),
    .X(\reg32_result.bit10.BitData ));
 sky130_fd_sc_hd__mux2_1 _0977_ (.A0(net3),
    .A1(net68),
    .S(_0448_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(_0457_),
    .X(\reg32_result.bit11.BitData ));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(net4),
    .A1(net161),
    .S(_0448_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0458_),
    .X(\reg32_result.bit12.BitData ));
 sky130_fd_sc_hd__buf_4 _0981_ (.A(\u1.q ),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(net5),
    .A1(net70),
    .S(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0460_),
    .X(\reg32_result.bit13.BitData ));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net6),
    .A1(net149),
    .S(_0459_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0461_),
    .X(\reg32_result.bit14.BitData ));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(net7),
    .A1(net147),
    .S(_0459_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(_0462_),
    .X(\reg32_result.bit15.BitData ));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(net8),
    .A1(net73),
    .S(_0459_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(_0463_),
    .X(\reg32_result.bit16.BitData ));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(net9),
    .A1(net74),
    .S(_0459_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(_0464_),
    .X(\reg32_result.bit17.BitData ));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(net10),
    .A1(net75),
    .S(_0459_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(_0465_),
    .X(\reg32_result.bit18.BitData ));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net11),
    .A1(net76),
    .S(_0459_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(_0466_),
    .X(\reg32_result.bit19.BitData ));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net13),
    .A1(net77),
    .S(_0459_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(_0467_),
    .X(\reg32_result.bit20.BitData ));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(net14),
    .A1(net79),
    .S(_0459_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(_0468_),
    .X(\reg32_result.bit21.BitData ));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(net15),
    .A1(net80),
    .S(_0459_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(_0469_),
    .X(\reg32_result.bit22.BitData ));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(net16),
    .A1(net81),
    .S(_0191_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0470_),
    .X(\reg32_result.bit23.BitData ));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(net17),
    .A1(net82),
    .S(_0191_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(_0471_),
    .X(\reg32_result.bit24.BitData ));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(net18),
    .A1(net83),
    .S(_0191_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(_0472_),
    .X(\reg32_result.bit25.BitData ));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(net19),
    .A1(net151),
    .S(_0191_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(_0473_),
    .X(\reg32_result.bit26.BitData ));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(net20),
    .A1(net85),
    .S(_0191_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(_0474_),
    .X(\reg32_result.bit27.BitData ));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(net21),
    .A1(net86),
    .S(_0191_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(_0475_),
    .X(\reg32_result.bit28.BitData ));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(net22),
    .A1(net140),
    .S(_0191_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(_0476_),
    .X(\reg32_result.bit29.BitData ));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(net24),
    .A1(net88),
    .S(_0191_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0477_),
    .X(\reg32_result.bit30.BitData ));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(net25),
    .A1(net90),
    .S(_0191_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(_0478_),
    .X(\reg32_result.bit31.BitData ));
 sky130_fd_sc_hd__or4_1 _1020_ (.A(net35),
    .B(net34),
    .C(net44),
    .D(net63),
    .X(_0479_));
 sky130_fd_sc_hd__or4_1 _1021_ (.A(net39),
    .B(net38),
    .C(net37),
    .D(net36),
    .X(_0480_));
 sky130_fd_sc_hd__or4_1 _1022_ (.A(net62),
    .B(net61),
    .C(net60),
    .D(net59),
    .X(_0481_));
 sky130_fd_sc_hd__or4_1 _1023_ (.A(net57),
    .B(net54),
    .C(net43),
    .D(net33),
    .X(_0482_));
 sky130_fd_sc_hd__or4_1 _1024_ (.A(_0479_),
    .B(_0480_),
    .C(_0481_),
    .D(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__or4_1 _1025_ (.A(net52),
    .B(net51),
    .C(net50),
    .D(net49),
    .X(_0484_));
 sky130_fd_sc_hd__or4_1 _1026_ (.A(net64),
    .B(net56),
    .C(net58),
    .D(net53),
    .X(_0485_));
 sky130_fd_sc_hd__or4_1 _1027_ (.A(net48),
    .B(net47),
    .C(net46),
    .D(net45),
    .X(_0486_));
 sky130_fd_sc_hd__or4_1 _1028_ (.A(net55),
    .B(net42),
    .C(net41),
    .D(net40),
    .X(_0487_));
 sky130_fd_sc_hd__or4_1 _1029_ (.A(_0484_),
    .B(_0485_),
    .C(_0486_),
    .D(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_1 _1030_ (.A(_0483_),
    .B(_0488_),
    .Y(net131));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(_0190_),
    .B(_0199_),
    .Y(\u1.d ));
 sky130_fd_sc_hd__buf_2 _1032_ (.A(net65),
    .X(_0489_));
 sky130_fd_sc_hd__buf_2 _1033_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__buf_2 _1034_ (.A(net66),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _1035_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and2b_1 _1036_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _1037_ (.A(_0493_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _1038_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(_0494_),
    .X(_0001_));
 sky130_fd_sc_hd__and2b_1 _1040_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(_0495_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _1042_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _1043_ (.A(_0496_),
    .X(_0003_));
 sky130_fd_sc_hd__and2b_1 _1044_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _1045_ (.A(_0497_),
    .X(_0004_));
 sky130_fd_sc_hd__and2b_1 _1046_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0498_),
    .X(_0005_));
 sky130_fd_sc_hd__and2b_1 _1048_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0499_),
    .X(_0006_));
 sky130_fd_sc_hd__and2b_1 _1050_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0500_),
    .X(_0007_));
 sky130_fd_sc_hd__and2b_1 _1052_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0501_),
    .X(_0008_));
 sky130_fd_sc_hd__and2b_1 _1054_ (.A_N(_0490_),
    .B(_0492_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0502_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _1056_ (.A(_0489_),
    .X(_0503_));
 sky130_fd_sc_hd__buf_2 _1057_ (.A(_0491_),
    .X(_0504_));
 sky130_fd_sc_hd__and2b_1 _1058_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1059_ (.A(_0505_),
    .X(_0010_));
 sky130_fd_sc_hd__and2b_1 _1060_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0506_),
    .X(_0011_));
 sky130_fd_sc_hd__and2b_1 _1062_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _1063_ (.A(_0507_),
    .X(_0012_));
 sky130_fd_sc_hd__and2b_1 _1064_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0508_),
    .X(_0013_));
 sky130_fd_sc_hd__and2b_1 _1066_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1067_ (.A(_0509_),
    .X(_0014_));
 sky130_fd_sc_hd__and2b_1 _1068_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _1069_ (.A(_0510_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _1070_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _1071_ (.A(_0511_),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _1072_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _1073_ (.A(_0512_),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _1074_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(_0513_),
    .X(_0018_));
 sky130_fd_sc_hd__and2b_1 _1076_ (.A_N(_0503_),
    .B(_0504_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _1077_ (.A(_0514_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_2 _1078_ (.A(_0489_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_2 _1079_ (.A(_0491_),
    .X(_0516_));
 sky130_fd_sc_hd__and2b_1 _1080_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1081_ (.A(_0517_),
    .X(_0020_));
 sky130_fd_sc_hd__and2b_1 _1082_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1083_ (.A(_0518_),
    .X(_0021_));
 sky130_fd_sc_hd__and2b_1 _1084_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _1085_ (.A(_0519_),
    .X(_0022_));
 sky130_fd_sc_hd__and2b_1 _1086_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _1087_ (.A(_0520_),
    .X(_0023_));
 sky130_fd_sc_hd__and2b_1 _1088_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0521_),
    .X(_0024_));
 sky130_fd_sc_hd__and2b_1 _1090_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _1091_ (.A(_0522_),
    .X(_0025_));
 sky130_fd_sc_hd__and2b_1 _1092_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _1093_ (.A(_0523_),
    .X(_0026_));
 sky130_fd_sc_hd__and2b_1 _1094_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _1095_ (.A(_0524_),
    .X(_0027_));
 sky130_fd_sc_hd__and2b_1 _1096_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _1097_ (.A(_0525_),
    .X(_0028_));
 sky130_fd_sc_hd__and2b_1 _1098_ (.A_N(_0515_),
    .B(_0516_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1099_ (.A(_0526_),
    .X(_0029_));
 sky130_fd_sc_hd__buf_2 _1100_ (.A(_0489_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _1101_ (.A(_0491_),
    .X(_0528_));
 sky130_fd_sc_hd__and2b_1 _1102_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _1103_ (.A(_0529_),
    .X(_0030_));
 sky130_fd_sc_hd__and2b_1 _1104_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1105_ (.A(_0530_),
    .X(_0031_));
 sky130_fd_sc_hd__and2b_1 _1106_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _1107_ (.A(_0531_),
    .X(_0032_));
 sky130_fd_sc_hd__and2b_1 _1108_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1109_ (.A(_0532_),
    .X(_0033_));
 sky130_fd_sc_hd__and2b_1 _1110_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_1 _1111_ (.A(_0533_),
    .X(_0034_));
 sky130_fd_sc_hd__and2b_1 _1112_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _1113_ (.A(_0534_),
    .X(_0035_));
 sky130_fd_sc_hd__and2b_1 _1114_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _1115_ (.A(_0535_),
    .X(_0036_));
 sky130_fd_sc_hd__and2b_1 _1116_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1117_ (.A(_0536_),
    .X(_0037_));
 sky130_fd_sc_hd__and2b_1 _1118_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _1119_ (.A(_0537_),
    .X(_0038_));
 sky130_fd_sc_hd__and2b_1 _1120_ (.A_N(_0527_),
    .B(_0528_),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1121_ (.A(_0538_),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_2 _1122_ (.A(_0489_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_2 _1123_ (.A(_0491_),
    .X(_0540_));
 sky130_fd_sc_hd__and2b_1 _1124_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _1125_ (.A(_0541_),
    .X(_0040_));
 sky130_fd_sc_hd__and2b_1 _1126_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _1127_ (.A(_0542_),
    .X(_0041_));
 sky130_fd_sc_hd__and2b_1 _1128_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1129_ (.A(_0543_),
    .X(_0042_));
 sky130_fd_sc_hd__and2b_1 _1130_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_1 _1131_ (.A(_0544_),
    .X(_0043_));
 sky130_fd_sc_hd__and2b_1 _1132_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0545_));
 sky130_fd_sc_hd__clkbuf_1 _1133_ (.A(_0545_),
    .X(_0044_));
 sky130_fd_sc_hd__and2b_1 _1134_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _1135_ (.A(_0546_),
    .X(_0045_));
 sky130_fd_sc_hd__and2b_1 _1136_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0547_));
 sky130_fd_sc_hd__clkbuf_1 _1137_ (.A(_0547_),
    .X(_0046_));
 sky130_fd_sc_hd__and2b_1 _1138_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _1139_ (.A(_0548_),
    .X(_0047_));
 sky130_fd_sc_hd__and2b_1 _1140_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0549_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0549_),
    .X(_0048_));
 sky130_fd_sc_hd__and2b_1 _1142_ (.A_N(_0539_),
    .B(_0540_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_1 _1143_ (.A(_0550_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_2 _1144_ (.A(_0489_),
    .X(_0551_));
 sky130_fd_sc_hd__buf_2 _1145_ (.A(_0491_),
    .X(_0552_));
 sky130_fd_sc_hd__and2b_1 _1146_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(_0553_),
    .X(_0050_));
 sky130_fd_sc_hd__and2b_1 _1148_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(_0554_),
    .X(_0051_));
 sky130_fd_sc_hd__and2b_1 _1150_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_1 _1151_ (.A(_0555_),
    .X(_0052_));
 sky130_fd_sc_hd__and2b_1 _1152_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0556_),
    .X(_0053_));
 sky130_fd_sc_hd__and2b_1 _1154_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _1155_ (.A(_0557_),
    .X(_0054_));
 sky130_fd_sc_hd__and2b_1 _1156_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_1 _1157_ (.A(_0558_),
    .X(_0055_));
 sky130_fd_sc_hd__and2b_1 _1158_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_1 _1159_ (.A(_0559_),
    .X(_0056_));
 sky130_fd_sc_hd__and2b_1 _1160_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _1161_ (.A(_0560_),
    .X(_0057_));
 sky130_fd_sc_hd__and2b_1 _1162_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _1163_ (.A(_0561_),
    .X(_0058_));
 sky130_fd_sc_hd__and2b_1 _1164_ (.A_N(_0551_),
    .B(_0552_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _1165_ (.A(_0562_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_2 _1166_ (.A(_0489_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_2 _1167_ (.A(_0491_),
    .X(_0564_));
 sky130_fd_sc_hd__and2b_1 _1168_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0565_),
    .X(_0060_));
 sky130_fd_sc_hd__and2b_1 _1170_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _1171_ (.A(_0566_),
    .X(_0061_));
 sky130_fd_sc_hd__and2b_1 _1172_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1173_ (.A(_0567_),
    .X(_0062_));
 sky130_fd_sc_hd__and2b_1 _1174_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_1 _1175_ (.A(_0568_),
    .X(_0063_));
 sky130_fd_sc_hd__and2b_1 _1176_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1177_ (.A(_0569_),
    .X(_0064_));
 sky130_fd_sc_hd__and2b_1 _1178_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _1179_ (.A(_0570_),
    .X(_0065_));
 sky130_fd_sc_hd__and2b_1 _1180_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0571_),
    .X(_0066_));
 sky130_fd_sc_hd__and2b_1 _1182_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _1183_ (.A(_0572_),
    .X(_0067_));
 sky130_fd_sc_hd__and2b_1 _1184_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_1 _1185_ (.A(_0573_),
    .X(_0068_));
 sky130_fd_sc_hd__and2b_1 _1186_ (.A_N(_0563_),
    .B(_0564_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _1187_ (.A(_0574_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_2 _1188_ (.A(_0489_),
    .X(_0575_));
 sky130_fd_sc_hd__buf_2 _1189_ (.A(_0491_),
    .X(_0576_));
 sky130_fd_sc_hd__and2b_1 _1190_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0577_),
    .X(_0070_));
 sky130_fd_sc_hd__and2b_1 _1192_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _1193_ (.A(_0578_),
    .X(_0071_));
 sky130_fd_sc_hd__and2b_1 _1194_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _1195_ (.A(_0579_),
    .X(_0072_));
 sky130_fd_sc_hd__and2b_1 _1196_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _1197_ (.A(_0580_),
    .X(_0073_));
 sky130_fd_sc_hd__and2b_1 _1198_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _1199_ (.A(_0581_),
    .X(_0074_));
 sky130_fd_sc_hd__and2b_1 _1200_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_1 _1201_ (.A(_0582_),
    .X(_0075_));
 sky130_fd_sc_hd__and2b_1 _1202_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _1203_ (.A(_0583_),
    .X(_0076_));
 sky130_fd_sc_hd__and2b_1 _1204_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0584_),
    .X(_0077_));
 sky130_fd_sc_hd__and2b_1 _1206_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _1207_ (.A(_0585_),
    .X(_0078_));
 sky130_fd_sc_hd__and2b_1 _1208_ (.A_N(_0575_),
    .B(_0576_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_1 _1209_ (.A(_0586_),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_2 _1210_ (.A(net65),
    .X(_0587_));
 sky130_fd_sc_hd__buf_2 _1211_ (.A(net66),
    .X(_0588_));
 sky130_fd_sc_hd__and2b_1 _1212_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__clkbuf_1 _1213_ (.A(_0589_),
    .X(_0080_));
 sky130_fd_sc_hd__and2b_1 _1214_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_1 _1215_ (.A(_0590_),
    .X(_0081_));
 sky130_fd_sc_hd__and2b_1 _1216_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_1 _1217_ (.A(_0591_),
    .X(_0082_));
 sky130_fd_sc_hd__and2b_1 _1218_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_1 _1219_ (.A(_0592_),
    .X(_0083_));
 sky130_fd_sc_hd__and2b_1 _1220_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _1221_ (.A(_0134_),
    .X(_0084_));
 sky130_fd_sc_hd__and2b_1 _1222_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _1223_ (.A(_0135_),
    .X(_0085_));
 sky130_fd_sc_hd__and2b_1 _1224_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1225_ (.A(_0136_),
    .X(_0086_));
 sky130_fd_sc_hd__and2b_1 _1226_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _1227_ (.A(_0137_),
    .X(_0087_));
 sky130_fd_sc_hd__and2b_1 _1228_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1229_ (.A(_0138_),
    .X(_0088_));
 sky130_fd_sc_hd__and2b_1 _1230_ (.A_N(_0587_),
    .B(_0588_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _1231_ (.A(_0139_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_2 _1232_ (.A(net65),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_2 _1233_ (.A(net66),
    .X(_0141_));
 sky130_fd_sc_hd__and2b_1 _1234_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _1235_ (.A(_0142_),
    .X(_0090_));
 sky130_fd_sc_hd__and2b_1 _1236_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _1237_ (.A(_0143_),
    .X(_0091_));
 sky130_fd_sc_hd__and2b_1 _1238_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _1239_ (.A(_0144_),
    .X(_0092_));
 sky130_fd_sc_hd__and2b_1 _1240_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _1241_ (.A(_0145_),
    .X(_0093_));
 sky130_fd_sc_hd__and2b_1 _1242_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _1243_ (.A(_0146_),
    .X(_0094_));
 sky130_fd_sc_hd__and2b_1 _1244_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _1245_ (.A(_0147_),
    .X(_0095_));
 sky130_fd_sc_hd__and2b_1 _1246_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _1247_ (.A(_0148_),
    .X(_0096_));
 sky130_fd_sc_hd__and2b_1 _1248_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _1249_ (.A(_0149_),
    .X(_0097_));
 sky130_fd_sc_hd__and2b_1 _1250_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _1251_ (.A(_0150_),
    .X(_0098_));
 sky130_fd_sc_hd__and2b_1 _1252_ (.A_N(_0140_),
    .B(_0141_),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _1253_ (.A(_0151_),
    .X(_0099_));
 sky130_fd_sc_hd__and2b_1 _1254_ (.A_N(_0489_),
    .B(_0491_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _1255_ (.A(_0152_),
    .X(_0100_));
 sky130_fd_sc_hd__and2b_1 _1256_ (.A_N(_0489_),
    .B(_0491_),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _1257_ (.A(_0153_),
    .X(_0101_));
 sky130_fd_sc_hd__dfrtp_4 _1258_ (.CLK(clknet_3_4__leaf_clk),
    .D(\u1.d ),
    .RESET_B(_0000_),
    .Q(\u1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(clknet_3_4__leaf_clk),
    .D(\cycle_reg.bit0.BitData ),
    .RESET_B(_0001_),
    .Q(\cycle_reg.bit0.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(clknet_3_4__leaf_clk),
    .D(\cycle_reg.bit1.BitData ),
    .RESET_B(_0002_),
    .Q(\cycle_reg.bit1.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(clknet_3_4__leaf_clk),
    .D(\cycle_reg.bit2.BitData ),
    .RESET_B(_0003_),
    .Q(\cycle_reg.bit2.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(clknet_3_4__leaf_clk),
    .D(\cycle_reg.bit3.BitData ),
    .RESET_B(_0004_),
    .Q(\cycle_reg.bit3.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(clknet_3_4__leaf_clk),
    .D(\cycle_reg.bit4.BitData ),
    .RESET_B(_0005_),
    .Q(\cycle_reg.bit4.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1264_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0102_),
    .RESET_B(_0006_),
    .Q(\reg32_denom.bit0.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0103_),
    .RESET_B(_0007_),
    .Q(\reg32_denom.bit19.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1266_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0104_),
    .RESET_B(_0008_),
    .Q(\reg32_denom.bit29.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1267_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0105_),
    .RESET_B(_0009_),
    .Q(\reg32_denom.bit31.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0106_),
    .RESET_B(_0010_),
    .Q(\reg32_denom.bit4.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1269_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0107_),
    .RESET_B(_0011_),
    .Q(\reg32_denom.bit5.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1270_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0108_),
    .RESET_B(_0012_),
    .Q(\reg32_denom.bit6.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1271_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0109_),
    .RESET_B(_0013_),
    .Q(\reg32_denom.bit7.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1272_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0110_),
    .RESET_B(_0014_),
    .Q(\reg32_denom.bit8.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1273_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0111_),
    .RESET_B(_0015_),
    .Q(\reg32_denom.bit1.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1274_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0112_),
    .RESET_B(_0016_),
    .Q(\reg32_denom.bit10.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1275_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0113_),
    .RESET_B(_0017_),
    .Q(\reg32_denom.bit11.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1276_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0114_),
    .RESET_B(_0018_),
    .Q(\reg32_denom.bit12.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1277_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0115_),
    .RESET_B(_0019_),
    .Q(\reg32_denom.bit13.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1278_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0116_),
    .RESET_B(_0020_),
    .Q(\reg32_denom.bit14.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1279_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0117_),
    .RESET_B(_0021_),
    .Q(\reg32_denom.bit15.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1280_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0118_),
    .RESET_B(_0022_),
    .Q(\reg32_denom.bit16.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1281_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0119_),
    .RESET_B(_0023_),
    .Q(\reg32_denom.bit17.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1282_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0120_),
    .RESET_B(_0024_),
    .Q(\reg32_denom.bit18.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1283_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0121_),
    .RESET_B(_0025_),
    .Q(\reg32_denom.bit2.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1284_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0122_),
    .RESET_B(_0026_),
    .Q(\reg32_denom.bit20.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1285_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0123_),
    .RESET_B(_0027_),
    .Q(\reg32_denom.bit21.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1286_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0124_),
    .RESET_B(_0028_),
    .Q(\reg32_denom.bit22.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1287_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0125_),
    .RESET_B(_0029_),
    .Q(\reg32_denom.bit23.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1288_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0126_),
    .RESET_B(_0030_),
    .Q(\reg32_denom.bit24.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1289_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0127_),
    .RESET_B(_0031_),
    .Q(\reg32_denom.bit25.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1290_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0128_),
    .RESET_B(_0032_),
    .Q(\reg32_denom.bit26.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1291_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0129_),
    .RESET_B(_0033_),
    .Q(\reg32_denom.bit27.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1292_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0130_),
    .RESET_B(_0034_),
    .Q(\reg32_denom.bit28.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1293_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0131_),
    .RESET_B(_0035_),
    .Q(\reg32_denom.bit3.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1294_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0132_),
    .RESET_B(_0036_),
    .Q(\reg32_denom.bit30.BitOut ));
 sky130_fd_sc_hd__dfrtp_1 _1295_ (.CLK(clknet_3_6__leaf_clk),
    .D(net158),
    .RESET_B(_0037_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_2 _1296_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_work.bit1.BitData ),
    .RESET_B(_0038_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_2 _1297_ (.CLK(clknet_3_4__leaf_clk),
    .D(\reg32_work.bit2.BitData ),
    .RESET_B(_0039_),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_2 _1298_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_work.bit3.BitData ),
    .RESET_B(_0040_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_2 _1299_ (.CLK(clknet_3_4__leaf_clk),
    .D(\reg32_work.bit4.BitData ),
    .RESET_B(_0041_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_2 _1300_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_work.bit5.BitData ),
    .RESET_B(_0042_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _1301_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_work.bit6.BitData ),
    .RESET_B(_0043_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_1 _1302_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_work.bit7.BitData ),
    .RESET_B(_0044_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_1 _1303_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_work.bit8.BitData ),
    .RESET_B(_0045_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_2 _1304_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_work.bit9.BitData ),
    .RESET_B(_0046_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_4 _1305_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_work.bit10.BitData ),
    .RESET_B(_0047_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _1306_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_work.bit11.BitData ),
    .RESET_B(_0048_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_2 _1307_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_work.bit12.BitData ),
    .RESET_B(_0049_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _1308_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_work.bit13.BitData ),
    .RESET_B(_0050_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _1309_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_work.bit14.BitData ),
    .RESET_B(_0051_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_2 _1310_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_work.bit15.BitData ),
    .RESET_B(_0052_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _1311_ (.CLK(clknet_3_1__leaf_clk),
    .D(\reg32_work.bit16.BitData ),
    .RESET_B(_0053_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _1312_ (.CLK(clknet_3_1__leaf_clk),
    .D(\reg32_work.bit17.BitData ),
    .RESET_B(_0054_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_2 _1313_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit18.BitData ),
    .RESET_B(_0055_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_2 _1314_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit19.BitData ),
    .RESET_B(_0056_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_2 _1315_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit20.BitData ),
    .RESET_B(_0057_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_2 _1316_ (.CLK(clknet_3_1__leaf_clk),
    .D(\reg32_work.bit21.BitData ),
    .RESET_B(_0058_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_2 _1317_ (.CLK(clknet_3_1__leaf_clk),
    .D(\reg32_work.bit22.BitData ),
    .RESET_B(_0059_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_1 _1318_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit23.BitData ),
    .RESET_B(_0060_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_2 _1319_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_work.bit24.BitData ),
    .RESET_B(_0061_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_2 _1320_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_work.bit25.BitData ),
    .RESET_B(_0062_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_2 _1321_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_work.bit26.BitData ),
    .RESET_B(_0063_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _1322_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_work.bit27.BitData ),
    .RESET_B(_0064_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_2 _1323_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_work.bit28.BitData ),
    .RESET_B(_0065_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_2 _1324_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_work.bit29.BitData ),
    .RESET_B(_0066_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_2 _1325_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit30.BitData ),
    .RESET_B(_0067_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_1 _1326_ (.CLK(clknet_3_0__leaf_clk),
    .D(\reg32_work.bit31.BitData ),
    .RESET_B(_0068_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_1 _1327_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0133_),
    .RESET_B(_0069_),
    .Q(\reg32_denom.bit9.BitOut ));
 sky130_fd_sc_hd__dfrtp_2 _1328_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit0.BitData ),
    .RESET_B(_0070_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _1329_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit1.BitData ),
    .RESET_B(_0071_),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _1330_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit2.BitData ),
    .RESET_B(_0072_),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _1331_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit3.BitData ),
    .RESET_B(_0073_),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _1332_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit4.BitData ),
    .RESET_B(_0074_),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _1333_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit5.BitData ),
    .RESET_B(_0075_),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _1334_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit6.BitData ),
    .RESET_B(_0076_),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_2 _1335_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit7.BitData ),
    .RESET_B(_0077_),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _1336_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit8.BitData ),
    .RESET_B(_0078_),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _1337_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit9.BitData ),
    .RESET_B(_0079_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _1338_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit10.BitData ),
    .RESET_B(_0080_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _1339_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit11.BitData ),
    .RESET_B(_0081_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _1340_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit12.BitData ),
    .RESET_B(_0082_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _1341_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_result.bit13.BitData ),
    .RESET_B(_0083_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1342_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_result.bit14.BitData ),
    .RESET_B(_0084_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _1343_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_result.bit15.BitData ),
    .RESET_B(_0085_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _1344_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit16.BitData ),
    .RESET_B(_0086_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _1345_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit17.BitData ),
    .RESET_B(_0087_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _1346_ (.CLK(clknet_3_7__leaf_clk),
    .D(\reg32_result.bit18.BitData ),
    .RESET_B(_0088_),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_4 _1347_ (.CLK(clknet_3_5__leaf_clk),
    .D(\reg32_result.bit19.BitData ),
    .RESET_B(_0089_),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _1348_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_result.bit20.BitData ),
    .RESET_B(_0090_),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_2 _1349_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_result.bit21.BitData ),
    .RESET_B(_0091_),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _1350_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit22.BitData ),
    .RESET_B(_0092_),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_2 _1351_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit23.BitData ),
    .RESET_B(_0093_),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _1352_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_result.bit24.BitData ),
    .RESET_B(_0094_),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _1353_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_result.bit25.BitData ),
    .RESET_B(_0095_),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _1354_ (.CLK(clknet_3_6__leaf_clk),
    .D(\reg32_result.bit26.BitData ),
    .RESET_B(_0096_),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_2 _1355_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit27.BitData ),
    .RESET_B(_0097_),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _1356_ (.CLK(clknet_3_2__leaf_clk),
    .D(\reg32_result.bit28.BitData ),
    .RESET_B(_0098_),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _1357_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit29.BitData ),
    .RESET_B(_0099_),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _1358_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit30.BitData ),
    .RESET_B(_0100_),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_2 _1359_ (.CLK(clknet_3_3__leaf_clk),
    .D(\reg32_result.bit31.BitData ),
    .RESET_B(_0101_),
    .Q(net91));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\cycle_reg.bit3.BitOut ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net106),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net129),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net120),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net114),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net72),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net110),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net71),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net121),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net84),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net89),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\cycle_reg.bit4.BitOut ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net105),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\reg32_denom.bit1.BitOut ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\reg32_denom.bit27.BitOut ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\reg32_denom.bit0.BitOut ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0331_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\reg32_work.bit0.BitData ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\reg32_denom.bit24.BitOut ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\reg32_denom.bit6.BitOut ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net69),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net108),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\cycle_reg.bit0.BitOut ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\reg32_denom.bit5.BitOut ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\reg32_denom.bit26.BitOut ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net78),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\reg32_denom.bit20.BitOut ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\cycle_reg.bit1.BitOut ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net118),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net124),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net87),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net128),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net111),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(reset),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(start),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap133 (.A(_0329_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(R[10]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(R[11]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(R[12]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(R[13]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(R[14]));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(R[15]));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(R[16]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(R[17]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(R[18]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(R[19]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(R[1]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(R[20]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(R[21]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(R[22]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(R[23]));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(R[24]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(R[25]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(R[26]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(R[27]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(R[28]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(R[29]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(R[2]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(R[30]));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net123),
    .X(R[31]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(R[3]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(R[4]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(R[5]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(R[6]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(R[7]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(R[8]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(R[9]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(err));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(ok));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(D[0]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(D[10]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(D[11]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(D[12]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(D[13]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(D[14]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(D[15]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(D[16]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(D[17]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(D[18]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(D[19]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(D[1]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(D[20]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(D[21]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(D[22]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(D[23]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(D[24]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(D[25]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(D[26]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(D[27]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(D[28]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(D[29]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(D[2]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(D[30]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(D[31]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(D[3]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(D[4]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(D[5]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(D[6]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(D[7]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(D[8]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(D[9]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(R[0]));
endmodule

