VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO divider
  CLASS BLOCK ;
  FOREIGN divider ;
  ORIGIN 0.000 0.000 ;
  SIZE 135.185 BY 145.905 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 115.640 135.185 116.240 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 141.905 77.650 145.905 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 3.440 135.185 4.040 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 132.640 135.185 133.240 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 141.905 87.310 145.905 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 141.905 16.470 145.905 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 40.840 135.185 41.440 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 108.840 135.185 109.440 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END A[21]
  PIN A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 141.905 129.170 145.905 ;
    END
  END A[22]
  PIN A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END A[23]
  PIN A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 112.240 135.185 112.840 ;
    END
  END A[24]
  PIN A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END A[25]
  PIN A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END A[26]
  PIN A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 54.440 135.185 55.040 ;
    END
  END A[27]
  PIN A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 0.040 135.185 0.640 ;
    END
  END A[28]
  PIN A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 17.040 135.185 17.640 ;
    END
  END A[29]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END A[2]
  PIN A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 141.905 29.350 145.905 ;
    END
  END A[30]
  PIN A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END A[31]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 141.905 109.850 145.905 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 91.840 135.185 92.440 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 141.905 45.450 145.905 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 141.905 26.130 145.905 ;
    END
  END B[0]
  PIN B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 141.905 116.290 145.905 ;
    END
  END B[10]
  PIN B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 81.640 135.185 82.240 ;
    END
  END B[11]
  PIN B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 85.040 135.185 85.640 ;
    END
  END B[12]
  PIN B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 141.905 61.550 145.905 ;
    END
  END B[13]
  PIN B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 141.905 64.770 145.905 ;
    END
  END B[14]
  PIN B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 141.905 48.670 145.905 ;
    END
  END B[15]
  PIN B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 141.905 90.530 145.905 ;
    END
  END B[16]
  PIN B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END B[17]
  PIN B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 141.905 3.590 145.905 ;
    END
  END B[18]
  PIN B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END B[19]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 61.240 135.185 61.840 ;
    END
  END B[1]
  PIN B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END B[20]
  PIN B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END B[21]
  PIN B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 37.440 135.185 38.040 ;
    END
  END B[22]
  PIN B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END B[23]
  PIN B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END B[24]
  PIN B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 141.905 13.250 145.905 ;
    END
  END B[25]
  PIN B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END B[26]
  PIN B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 141.905 122.730 145.905 ;
    END
  END B[27]
  PIN B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END B[28]
  PIN B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 142.840 135.185 143.440 ;
    END
  END B[29]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END B[2]
  PIN B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 102.040 135.185 102.640 ;
    END
  END B[30]
  PIN B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END B[31]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 141.905 132.390 145.905 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 141.905 32.570 145.905 ;
    END
  END B[9]
  PIN D[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.930 141.905 71.210 145.905 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 141.905 106.630 145.905 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 141.905 10.030 145.905 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 141.905 42.230 145.905 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 141.905 55.110 145.905 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 64.640 135.185 65.240 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 131.185 47.640 135.185 48.240 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 131.185 129.240 135.185 129.840 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 6.840 135.185 7.440 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 51.040 135.185 51.640 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 30.640 135.185 31.240 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 71.440 135.185 72.040 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 131.185 139.440 135.185 140.040 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 20.440 135.185 21.040 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 141.905 58.330 145.905 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 131.185 13.640 135.185 14.240 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 98.640 135.185 99.240 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END D[9]
  PIN R[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 131.185 34.040 135.185 34.640 ;
    END
  END R[0]
  PIN R[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END R[10]
  PIN R[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 78.240 135.185 78.840 ;
    END
  END R[11]
  PIN R[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 119.040 135.185 119.640 ;
    END
  END R[12]
  PIN R[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END R[13]
  PIN R[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 125.840 135.185 126.440 ;
    END
  END R[14]
  PIN R[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END R[15]
  PIN R[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END R[16]
  PIN R[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END R[17]
  PIN R[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END R[18]
  PIN R[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END R[19]
  PIN R[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END R[1]
  PIN R[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 141.905 35.790 145.905 ;
    END
  END R[20]
  PIN R[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 141.905 84.090 145.905 ;
    END
  END R[21]
  PIN R[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END R[22]
  PIN R[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END R[23]
  PIN R[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END R[24]
  PIN R[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.130 141.905 103.410 145.905 ;
    END
  END R[25]
  PIN R[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 141.905 74.430 145.905 ;
    END
  END R[26]
  PIN R[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END R[27]
  PIN R[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.230 141.905 119.510 145.905 ;
    END
  END R[28]
  PIN R[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 23.840 135.185 24.440 ;
    END
  END R[29]
  PIN R[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END R[2]
  PIN R[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END R[30]
  PIN R[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END R[31]
  PIN R[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END R[3]
  PIN R[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END R[4]
  PIN R[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 95.240 135.185 95.840 ;
    END
  END R[5]
  PIN R[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END R[6]
  PIN R[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 99.910 141.905 100.190 145.905 ;
    END
  END R[7]
  PIN R[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 141.905 93.750 145.905 ;
    END
  END R[8]
  PIN R[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 141.905 0.370 145.905 ;
    END
  END R[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.485 10.640 25.085 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.420 10.640 56.020 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.355 10.640 86.955 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.290 10.640 117.890 133.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 28.680 129.500 30.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 59.280 129.500 60.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 89.880 129.500 91.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 120.480 129.500 122.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.185 10.640 21.785 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.120 10.640 52.720 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.055 10.640 83.655 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.990 10.640 114.590 133.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 25.380 129.500 26.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 55.980 129.500 57.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 86.580 129.500 88.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 117.180 129.500 118.780 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 141.905 19.690 145.905 ;
    END
  END clk
  PIN err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END err
  PIN ok
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END ok
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END reset
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 131.185 68.040 135.185 68.640 ;
    END
  END start
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 129.260 133.365 ;
      LAYER met1 ;
        RECT 0.070 7.520 132.410 133.520 ;
      LAYER met2 ;
        RECT 0.650 141.625 3.030 143.325 ;
        RECT 3.870 141.625 9.470 143.325 ;
        RECT 10.310 141.625 12.690 143.325 ;
        RECT 13.530 141.625 15.910 143.325 ;
        RECT 16.750 141.625 19.130 143.325 ;
        RECT 19.970 141.625 25.570 143.325 ;
        RECT 26.410 141.625 28.790 143.325 ;
        RECT 29.630 141.625 32.010 143.325 ;
        RECT 32.850 141.625 35.230 143.325 ;
        RECT 36.070 141.625 41.670 143.325 ;
        RECT 42.510 141.625 44.890 143.325 ;
        RECT 45.730 141.625 48.110 143.325 ;
        RECT 48.950 141.625 54.550 143.325 ;
        RECT 55.390 141.625 57.770 143.325 ;
        RECT 58.610 141.625 60.990 143.325 ;
        RECT 61.830 141.625 64.210 143.325 ;
        RECT 65.050 141.625 70.650 143.325 ;
        RECT 71.490 141.625 73.870 143.325 ;
        RECT 74.710 141.625 77.090 143.325 ;
        RECT 77.930 141.625 83.530 143.325 ;
        RECT 84.370 141.625 86.750 143.325 ;
        RECT 87.590 141.625 89.970 143.325 ;
        RECT 90.810 141.625 93.190 143.325 ;
        RECT 94.030 141.625 99.630 143.325 ;
        RECT 100.470 141.625 102.850 143.325 ;
        RECT 103.690 141.625 106.070 143.325 ;
        RECT 106.910 141.625 109.290 143.325 ;
        RECT 110.130 141.625 115.730 143.325 ;
        RECT 116.570 141.625 118.950 143.325 ;
        RECT 119.790 141.625 122.170 143.325 ;
        RECT 123.010 141.625 128.610 143.325 ;
        RECT 129.450 141.625 131.830 143.325 ;
        RECT 0.100 4.280 132.380 141.625 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 132.380 4.280 ;
      LAYER met3 ;
        RECT 4.400 142.440 130.785 143.305 ;
        RECT 3.990 140.440 131.955 142.440 ;
        RECT 3.990 139.040 130.785 140.440 ;
        RECT 3.990 137.040 131.955 139.040 ;
        RECT 4.400 135.640 131.955 137.040 ;
        RECT 3.990 133.640 131.955 135.640 ;
        RECT 4.400 132.240 130.785 133.640 ;
        RECT 3.990 130.240 131.955 132.240 ;
        RECT 4.400 128.840 130.785 130.240 ;
        RECT 3.990 126.840 131.955 128.840 ;
        RECT 4.400 125.440 130.785 126.840 ;
        RECT 3.990 120.040 131.955 125.440 ;
        RECT 4.400 118.640 130.785 120.040 ;
        RECT 3.990 116.640 131.955 118.640 ;
        RECT 4.400 115.240 130.785 116.640 ;
        RECT 3.990 113.240 131.955 115.240 ;
        RECT 4.400 111.840 130.785 113.240 ;
        RECT 3.990 109.840 131.955 111.840 ;
        RECT 3.990 108.440 130.785 109.840 ;
        RECT 3.990 106.440 131.955 108.440 ;
        RECT 4.400 105.040 131.955 106.440 ;
        RECT 3.990 103.040 131.955 105.040 ;
        RECT 4.400 101.640 130.785 103.040 ;
        RECT 3.990 99.640 131.955 101.640 ;
        RECT 4.400 98.240 130.785 99.640 ;
        RECT 3.990 96.240 131.955 98.240 ;
        RECT 4.400 94.840 130.785 96.240 ;
        RECT 3.990 92.840 131.955 94.840 ;
        RECT 3.990 91.440 130.785 92.840 ;
        RECT 3.990 89.440 131.955 91.440 ;
        RECT 4.400 88.040 131.955 89.440 ;
        RECT 3.990 86.040 131.955 88.040 ;
        RECT 4.400 84.640 130.785 86.040 ;
        RECT 3.990 82.640 131.955 84.640 ;
        RECT 4.400 81.240 130.785 82.640 ;
        RECT 3.990 79.240 131.955 81.240 ;
        RECT 4.400 77.840 130.785 79.240 ;
        RECT 3.990 72.440 131.955 77.840 ;
        RECT 4.400 71.040 130.785 72.440 ;
        RECT 3.990 69.040 131.955 71.040 ;
        RECT 4.400 67.640 130.785 69.040 ;
        RECT 3.990 65.640 131.955 67.640 ;
        RECT 4.400 64.240 130.785 65.640 ;
        RECT 3.990 62.240 131.955 64.240 ;
        RECT 3.990 60.840 130.785 62.240 ;
        RECT 3.990 58.840 131.955 60.840 ;
        RECT 4.400 57.440 131.955 58.840 ;
        RECT 3.990 55.440 131.955 57.440 ;
        RECT 4.400 54.040 130.785 55.440 ;
        RECT 3.990 52.040 131.955 54.040 ;
        RECT 4.400 50.640 130.785 52.040 ;
        RECT 3.990 48.640 131.955 50.640 ;
        RECT 4.400 47.240 130.785 48.640 ;
        RECT 3.990 41.840 131.955 47.240 ;
        RECT 4.400 40.440 130.785 41.840 ;
        RECT 3.990 38.440 131.955 40.440 ;
        RECT 4.400 37.040 130.785 38.440 ;
        RECT 3.990 35.040 131.955 37.040 ;
        RECT 4.400 33.640 130.785 35.040 ;
        RECT 3.990 31.640 131.955 33.640 ;
        RECT 3.990 30.240 130.785 31.640 ;
        RECT 3.990 28.240 131.955 30.240 ;
        RECT 4.400 26.840 131.955 28.240 ;
        RECT 3.990 24.840 131.955 26.840 ;
        RECT 4.400 23.440 130.785 24.840 ;
        RECT 3.990 21.440 131.955 23.440 ;
        RECT 4.400 20.040 130.785 21.440 ;
        RECT 3.990 18.040 131.955 20.040 ;
        RECT 4.400 16.640 130.785 18.040 ;
        RECT 3.990 14.640 131.955 16.640 ;
        RECT 3.990 13.240 130.785 14.640 ;
        RECT 3.990 11.240 131.955 13.240 ;
        RECT 4.400 9.840 131.955 11.240 ;
        RECT 3.990 7.840 131.955 9.840 ;
        RECT 4.400 6.440 130.785 7.840 ;
        RECT 3.990 4.440 131.955 6.440 ;
        RECT 4.400 3.040 130.785 4.440 ;
        RECT 3.990 1.040 131.955 3.040 ;
        RECT 3.990 0.175 130.785 1.040 ;
      LAYER met4 ;
        RECT 38.935 13.095 50.720 123.585 ;
        RECT 53.120 13.095 54.020 123.585 ;
        RECT 56.420 13.095 76.985 123.585 ;
  END
END divider
END LIBRARY

